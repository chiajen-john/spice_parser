*
*
*
*                       LINUX           Thu Nov 23 19:11:37 2023
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 19.1.3-s062
*  Build Date     : Tue Jul 23 02:42:20 PDT 2019
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT bit_cell_col_64 VDD VSS WL<0> WL<10> WL<11> WL<12> WL<13> WL<14> WL<15>
+ WL<16> WL<17> WL<18> WL<19> WL<1> WL<20> WL<21> WL<22> WL<23> WL<24> WL<25>
+ WL<26> WL<27> WL<28> WL<29> WL<2> WL<30> WL<31> WL<32> WL<33> WL<34> WL<35>
+ WL<36> WL<37> WL<38> WL<39> WL<3> WL<40> WL<41> WL<42> WL<43> WL<44> WL<45>
+ WL<46> WL<47> WL<48> WL<49> WL<4> WL<50> WL<51> WL<52> WL<53> WL<54> WL<55>
+ WL<56> WL<57> WL<58> WL<59> WL<5> WL<60> WL<61> WL<62> WL<63> WL<6> WL<7>
+ WL<8> WL<9> BL BLB
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MI0<3>/I0<3>/I0<3>/NM0	I0<3>/I0<3>/I0<3>/Q#6	WL<63>#1	BL#1	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<3>/NM2	I0<3>/I0<3>/I0<3>/Q#6	I0<3>/I0<3>/I0<3>/QB#3	VSS#4
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I0<3>/I0<3>/NM1	BLB#1	WL<63>#3	I0<3>/I0<3>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I0<3>/I0<3>/NM3	I0<3>/I0<3>/I0<3>/QB#4	I0<3>/I0<3>/I0<3>/Q	VSS#73
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<1>/NM0	I0<3>/I0<3>/I0<1>/Q#6	WL<61>#1	BL#3	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<1>/NM2	I0<3>/I0<3>/I0<1>/Q#6	I0<3>/I0<3>/I0<1>/QB#3	VSS#6
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<1>/NM1	BLB#3	WL<61>#3	I0<3>/I0<3>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<1>/NM3	I0<3>/I0<3>/I0<1>/QB#4	I0<3>/I0<3>/I0<1>/Q	VSS#75
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<2>/NM0	I0<3>/I0<3>/I0<2>/Q#6	WL<62>#1	BL#1	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<2>/NM2	I0<3>/I0<3>/I0<2>/Q#6	I0<3>/I0<3>/I0<2>/QB#2	VSS#6
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<2>/NM1	BLB#3	WL<62>#4	I0<3>/I0<3>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<2>/NM3	I0<3>/I0<3>/I0<2>/QB#4	I0<3>/I0<3>/I0<2>/Q	VSS#73
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<0>/NM0	I0<3>/I0<3>/I0<0>/Q#6	WL<60>#1	BL#3	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<0>/NM2	I0<3>/I0<3>/I0<0>/Q#6	I0<3>/I0<3>/I0<0>/QB#2	VSS#8
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<0>/NM1	BLB#5	WL<60>#4	I0<3>/I0<3>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<3>/I0<0>/NM3	I0<3>/I0<3>/I0<0>/QB#4	I0<3>/I0<3>/I0<0>/Q	VSS#75
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<3>/NM0	I0<3>/I0<2>/I0<3>/Q#6	WL<59>#1	BL#5	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<3>/NM2	I0<3>/I0<2>/I0<3>/Q#6	I0<3>/I0<2>/I0<3>/QB#3	VSS#8
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<3>/NM1	BLB#5	WL<59>#3	I0<3>/I0<2>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<3>/NM3	I0<3>/I0<2>/I0<3>/QB#4	I0<3>/I0<2>/I0<3>/Q	VSS#77
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<1>/NM0	I0<3>/I0<2>/I0<1>/Q#6	WL<57>#1	BL#7	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<1>/NM2	I0<3>/I0<2>/I0<1>/Q#6	I0<3>/I0<2>/I0<1>/QB#3	VSS#10
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<1>/NM1	BLB#7	WL<57>#3	I0<3>/I0<2>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<1>/NM3	I0<3>/I0<2>/I0<1>/QB#4	I0<3>/I0<2>/I0<1>/Q	VSS#79
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<2>/NM0	I0<3>/I0<2>/I0<2>/Q#6	WL<58>#1	BL#5	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<2>/NM2	I0<3>/I0<2>/I0<2>/Q#6	I0<3>/I0<2>/I0<2>/QB#2	VSS#10
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<2>/NM1	BLB#7	WL<58>#4	I0<3>/I0<2>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<2>/NM3	I0<3>/I0<2>/I0<2>/QB#4	I0<3>/I0<2>/I0<2>/Q	VSS#77
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<0>/NM0	I0<3>/I0<2>/I0<0>/Q#6	WL<56>#1	BL#7	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<0>/NM2	I0<3>/I0<2>/I0<0>/Q#6	I0<3>/I0<2>/I0<0>/QB#2	VSS#12
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<2>/I0<0>/NM1	BLB#9	WL<56>#4	I0<3>/I0<2>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<2>/I0<0>/NM3	I0<3>/I0<2>/I0<0>/QB#4	I0<3>/I0<2>/I0<0>/Q	VSS#79
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<3>/NM0	I0<3>/I0<1>/I0<3>/Q#6	WL<55>#1	BL#9	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<3>/NM2	I0<3>/I0<1>/I0<3>/Q#6	I0<3>/I0<1>/I0<3>/QB#3	VSS#12
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<3>/NM1	BLB#9	WL<55>#3	I0<3>/I0<1>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<3>/NM3	I0<3>/I0<1>/I0<3>/QB#4	I0<3>/I0<1>/I0<3>/Q	VSS#81
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<1>/NM0	I0<3>/I0<1>/I0<1>/Q#6	WL<53>#1	BL#11	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<1>/NM2	I0<3>/I0<1>/I0<1>/Q#6	I0<3>/I0<1>/I0<1>/QB#3	VSS#14
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<1>/NM1	BLB#11	WL<53>#3	I0<3>/I0<1>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<1>/NM3	I0<3>/I0<1>/I0<1>/QB#4	I0<3>/I0<1>/I0<1>/Q	VSS#83
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<2>/NM0	I0<3>/I0<1>/I0<2>/Q#6	WL<54>#1	BL#9	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<2>/NM2	I0<3>/I0<1>/I0<2>/Q#6	I0<3>/I0<1>/I0<2>/QB#2	VSS#14
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<2>/NM1	BLB#11	WL<54>#4	I0<3>/I0<1>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<2>/NM3	I0<3>/I0<1>/I0<2>/QB#4	I0<3>/I0<1>/I0<2>/Q	VSS#81
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<0>/NM0	I0<3>/I0<1>/I0<0>/Q#6	WL<52>#1	BL#11	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<0>/NM2	I0<3>/I0<1>/I0<0>/Q#6	I0<3>/I0<1>/I0<0>/QB#2	VSS#16
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<1>/I0<0>/NM1	BLB#13	WL<52>#4	I0<3>/I0<1>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<1>/I0<0>/NM3	I0<3>/I0<1>/I0<0>/QB#4	I0<3>/I0<1>/I0<0>/Q	VSS#83
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<3>/NM0	I0<3>/I0<0>/I0<3>/Q#6	WL<51>#1	BL#13	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<3>/NM2	I0<3>/I0<0>/I0<3>/Q#6	I0<3>/I0<0>/I0<3>/QB#3	VSS#16
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<3>/NM1	BLB#13	WL<51>#3	I0<3>/I0<0>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<3>/NM3	I0<3>/I0<0>/I0<3>/QB#4	I0<3>/I0<0>/I0<3>/Q	VSS#85
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<1>/NM0	I0<3>/I0<0>/I0<1>/Q#6	WL<49>#1	BL#15	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<1>/NM2	I0<3>/I0<0>/I0<1>/Q#6	I0<3>/I0<0>/I0<1>/QB#3	VSS#18
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<1>/NM1	BLB#15	WL<49>#3	I0<3>/I0<0>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<1>/NM3	I0<3>/I0<0>/I0<1>/QB#4	I0<3>/I0<0>/I0<1>/Q	VSS#87
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<2>/NM0	I0<3>/I0<0>/I0<2>/Q#6	WL<50>#1	BL#13	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<2>/NM2	I0<3>/I0<0>/I0<2>/Q#6	I0<3>/I0<0>/I0<2>/QB#2	VSS#18
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<2>/NM1	BLB#15	WL<50>#4	I0<3>/I0<0>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<2>/NM3	I0<3>/I0<0>/I0<2>/QB#4	I0<3>/I0<0>/I0<2>/Q	VSS#85
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<0>/NM0	I0<3>/I0<0>/I0<0>/Q#6	WL<48>#1	BL#15	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<0>/NM2	I0<3>/I0<0>/I0<0>/Q#6	I0<3>/I0<0>/I0<0>/QB#2	VSS#20
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<0>/I0<0>/NM1	BLB#17	WL<48>#4	I0<3>/I0<0>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<3>/I0<0>/I0<0>/NM3	I0<3>/I0<0>/I0<0>/QB#4	I0<3>/I0<0>/I0<0>/Q	VSS#87
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<3>/NM0	I0<2>/I0<3>/I0<3>/Q#6	WL<47>#1	BL#17	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<3>/NM2	I0<2>/I0<3>/I0<3>/Q#6	I0<2>/I0<3>/I0<3>/QB#3	VSS#20
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<3>/NM1	BLB#17	WL<47>#3	I0<2>/I0<3>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<3>/NM3	I0<2>/I0<3>/I0<3>/QB#4	I0<2>/I0<3>/I0<3>/Q	VSS#89
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<1>/NM0	I0<2>/I0<3>/I0<1>/Q#6	WL<45>#1	BL#19	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<1>/NM2	I0<2>/I0<3>/I0<1>/Q#6	I0<2>/I0<3>/I0<1>/QB#3	VSS#22
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<1>/NM1	BLB#19	WL<45>#3	I0<2>/I0<3>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<1>/NM3	I0<2>/I0<3>/I0<1>/QB#4	I0<2>/I0<3>/I0<1>/Q	VSS#91
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<2>/NM0	I0<2>/I0<3>/I0<2>/Q#6	WL<46>#1	BL#17	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<2>/NM2	I0<2>/I0<3>/I0<2>/Q#6	I0<2>/I0<3>/I0<2>/QB#2	VSS#22
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<2>/NM1	BLB#19	WL<46>#4	I0<2>/I0<3>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<2>/NM3	I0<2>/I0<3>/I0<2>/QB#4	I0<2>/I0<3>/I0<2>/Q	VSS#89
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<0>/NM0	I0<2>/I0<3>/I0<0>/Q#6	WL<44>#1	BL#19	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<0>/NM2	I0<2>/I0<3>/I0<0>/Q#6	I0<2>/I0<3>/I0<0>/QB#2	VSS#24
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<3>/I0<0>/NM1	BLB#21	WL<44>#4	I0<2>/I0<3>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<3>/I0<0>/NM3	I0<2>/I0<3>/I0<0>/QB#4	I0<2>/I0<3>/I0<0>/Q	VSS#91
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<3>/NM0	I0<2>/I0<2>/I0<3>/Q#6	WL<43>#1	BL#21	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<3>/NM2	I0<2>/I0<2>/I0<3>/Q#6	I0<2>/I0<2>/I0<3>/QB#3	VSS#24
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<3>/NM1	BLB#21	WL<43>#3	I0<2>/I0<2>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<3>/NM3	I0<2>/I0<2>/I0<3>/QB#4	I0<2>/I0<2>/I0<3>/Q	VSS#93
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<1>/NM0	I0<2>/I0<2>/I0<1>/Q#6	WL<41>#1	BL#23	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<1>/NM2	I0<2>/I0<2>/I0<1>/Q#6	I0<2>/I0<2>/I0<1>/QB#3	VSS#26
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<1>/NM1	BLB#23	WL<41>#3	I0<2>/I0<2>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<1>/NM3	I0<2>/I0<2>/I0<1>/QB#4	I0<2>/I0<2>/I0<1>/Q	VSS#95
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<2>/NM0	I0<2>/I0<2>/I0<2>/Q#6	WL<42>#1	BL#21	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<2>/NM2	I0<2>/I0<2>/I0<2>/Q#6	I0<2>/I0<2>/I0<2>/QB#2	VSS#26
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<2>/NM1	BLB#23	WL<42>#4	I0<2>/I0<2>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<2>/NM3	I0<2>/I0<2>/I0<2>/QB#4	I0<2>/I0<2>/I0<2>/Q	VSS#93
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<0>/NM0	I0<2>/I0<2>/I0<0>/Q#6	WL<40>#1	BL#23	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<0>/NM2	I0<2>/I0<2>/I0<0>/Q#6	I0<2>/I0<2>/I0<0>/QB#2	VSS#28
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<2>/I0<0>/NM1	BLB#25	WL<40>#4	I0<2>/I0<2>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<2>/I0<0>/NM3	I0<2>/I0<2>/I0<0>/QB#4	I0<2>/I0<2>/I0<0>/Q	VSS#95
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<3>/NM0	I0<2>/I0<1>/I0<3>/Q#6	WL<39>#1	BL#25	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<3>/NM2	I0<2>/I0<1>/I0<3>/Q#6	I0<2>/I0<1>/I0<3>/QB#3	VSS#28
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<3>/NM1	BLB#25	WL<39>#3	I0<2>/I0<1>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<3>/NM3	I0<2>/I0<1>/I0<3>/QB#4	I0<2>/I0<1>/I0<3>/Q	VSS#97
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<1>/NM0	I0<2>/I0<1>/I0<1>/Q#6	WL<37>#1	BL#27	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<1>/NM2	I0<2>/I0<1>/I0<1>/Q#6	I0<2>/I0<1>/I0<1>/QB#3	VSS#30
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<1>/NM1	BLB#27	WL<37>#3	I0<2>/I0<1>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<1>/NM3	I0<2>/I0<1>/I0<1>/QB#4	I0<2>/I0<1>/I0<1>/Q	VSS#99
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<2>/NM0	I0<2>/I0<1>/I0<2>/Q#6	WL<38>#1	BL#25	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<2>/NM2	I0<2>/I0<1>/I0<2>/Q#6	I0<2>/I0<1>/I0<2>/QB#2	VSS#30
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<2>/NM1	BLB#27	WL<38>#4	I0<2>/I0<1>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<2>/NM3	I0<2>/I0<1>/I0<2>/QB#4	I0<2>/I0<1>/I0<2>/Q	VSS#97
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<0>/NM0	I0<2>/I0<1>/I0<0>/Q#6	WL<36>#1	BL#27	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<0>/NM2	I0<2>/I0<1>/I0<0>/Q#6	I0<2>/I0<1>/I0<0>/QB#2	VSS#32
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<1>/I0<0>/NM1	BLB#29	WL<36>#4	I0<2>/I0<1>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<1>/I0<0>/NM3	I0<2>/I0<1>/I0<0>/QB#4	I0<2>/I0<1>/I0<0>/Q	VSS#99
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<3>/NM0	I0<2>/I0<0>/I0<3>/Q#6	WL<35>#1	BL#29	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<3>/NM2	I0<2>/I0<0>/I0<3>/Q#6	I0<2>/I0<0>/I0<3>/QB#3	VSS#32
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<3>/NM1	BLB#29	WL<35>#3	I0<2>/I0<0>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<3>/NM3	I0<2>/I0<0>/I0<3>/QB#4	I0<2>/I0<0>/I0<3>/Q	VSS#101
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<1>/NM0	I0<2>/I0<0>/I0<1>/Q#6	WL<33>#1	BL#31	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<1>/NM2	I0<2>/I0<0>/I0<1>/Q#6	I0<2>/I0<0>/I0<1>/QB#3	VSS#34
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<1>/NM1	BLB#31	WL<33>#3	I0<2>/I0<0>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<1>/NM3	I0<2>/I0<0>/I0<1>/QB#4	I0<2>/I0<0>/I0<1>/Q	VSS#103
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<2>/NM0	I0<2>/I0<0>/I0<2>/Q#6	WL<34>#1	BL#29	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<2>/NM2	I0<2>/I0<0>/I0<2>/Q#6	I0<2>/I0<0>/I0<2>/QB#2	VSS#34
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<2>/NM1	BLB#31	WL<34>#4	I0<2>/I0<0>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<2>/NM3	I0<2>/I0<0>/I0<2>/QB#4	I0<2>/I0<0>/I0<2>/Q	VSS#101
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<0>/NM0	I0<2>/I0<0>/I0<0>/Q#6	WL<32>#1	BL#31	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<0>/NM2	I0<2>/I0<0>/I0<0>/Q#6	I0<2>/I0<0>/I0<0>/QB#2	VSS#36
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<2>/I0<0>/I0<0>/NM1	BLB#33	WL<32>#4	I0<2>/I0<0>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<2>/I0<0>/I0<0>/NM3	I0<2>/I0<0>/I0<0>/QB#4	I0<2>/I0<0>/I0<0>/Q	VSS#103
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<3>/NM0	I0<1>/I0<3>/I0<3>/Q#6	WL<31>#1	BL#33	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<3>/NM2	I0<1>/I0<3>/I0<3>/Q#6	I0<1>/I0<3>/I0<3>/QB#3	VSS#36
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<3>/NM1	BLB#33	WL<31>#3	I0<1>/I0<3>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<3>/NM3	I0<1>/I0<3>/I0<3>/QB#4	I0<1>/I0<3>/I0<3>/Q	VSS#105
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<1>/NM0	I0<1>/I0<3>/I0<1>/Q#6	WL<29>#1	BL#35	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<1>/NM2	I0<1>/I0<3>/I0<1>/Q#6	I0<1>/I0<3>/I0<1>/QB#3	VSS#38
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<1>/NM1	BLB#35	WL<29>#3	I0<1>/I0<3>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<1>/NM3	I0<1>/I0<3>/I0<1>/QB#4	I0<1>/I0<3>/I0<1>/Q	VSS#107
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<2>/NM0	I0<1>/I0<3>/I0<2>/Q#6	WL<30>#1	BL#33	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<2>/NM2	I0<1>/I0<3>/I0<2>/Q#6	I0<1>/I0<3>/I0<2>/QB#2	VSS#38
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<2>/NM1	BLB#35	WL<30>#4	I0<1>/I0<3>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<2>/NM3	I0<1>/I0<3>/I0<2>/QB#4	I0<1>/I0<3>/I0<2>/Q	VSS#105
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<0>/NM0	I0<1>/I0<3>/I0<0>/Q#6	WL<28>#1	BL#35	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<0>/NM2	I0<1>/I0<3>/I0<0>/Q#6	I0<1>/I0<3>/I0<0>/QB#2	VSS#40
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<3>/I0<0>/NM1	BLB#37	WL<28>#4	I0<1>/I0<3>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<3>/I0<0>/NM3	I0<1>/I0<3>/I0<0>/QB#4	I0<1>/I0<3>/I0<0>/Q	VSS#107
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<3>/NM0	I0<1>/I0<2>/I0<3>/Q#6	WL<27>#1	BL#37	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<3>/NM2	I0<1>/I0<2>/I0<3>/Q#6	I0<1>/I0<2>/I0<3>/QB#3	VSS#40
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<3>/NM1	BLB#37	WL<27>#3	I0<1>/I0<2>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<3>/NM3	I0<1>/I0<2>/I0<3>/QB#4	I0<1>/I0<2>/I0<3>/Q	VSS#109
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<1>/NM0	I0<1>/I0<2>/I0<1>/Q#6	WL<25>#1	BL#39	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<1>/NM2	I0<1>/I0<2>/I0<1>/Q#6	I0<1>/I0<2>/I0<1>/QB#3	VSS#42
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<1>/NM1	BLB#39	WL<25>#3	I0<1>/I0<2>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<1>/NM3	I0<1>/I0<2>/I0<1>/QB#4	I0<1>/I0<2>/I0<1>/Q	VSS#111
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<2>/NM0	I0<1>/I0<2>/I0<2>/Q#6	WL<26>#1	BL#37	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<2>/NM2	I0<1>/I0<2>/I0<2>/Q#6	I0<1>/I0<2>/I0<2>/QB#2	VSS#42
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<2>/NM1	BLB#39	WL<26>#4	I0<1>/I0<2>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<2>/NM3	I0<1>/I0<2>/I0<2>/QB#4	I0<1>/I0<2>/I0<2>/Q	VSS#109
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<0>/NM0	I0<1>/I0<2>/I0<0>/Q#6	WL<24>#1	BL#39	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<0>/NM2	I0<1>/I0<2>/I0<0>/Q#6	I0<1>/I0<2>/I0<0>/QB#2	VSS#44
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<2>/I0<0>/NM1	BLB#41	WL<24>#4	I0<1>/I0<2>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<2>/I0<0>/NM3	I0<1>/I0<2>/I0<0>/QB#4	I0<1>/I0<2>/I0<0>/Q	VSS#111
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<3>/NM0	I0<1>/I0<1>/I0<3>/Q#6	WL<23>#1	BL#41	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<3>/NM2	I0<1>/I0<1>/I0<3>/Q#6	I0<1>/I0<1>/I0<3>/QB#3	VSS#44
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<3>/NM1	BLB#41	WL<23>#3	I0<1>/I0<1>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<3>/NM3	I0<1>/I0<1>/I0<3>/QB#4	I0<1>/I0<1>/I0<3>/Q	VSS#113
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<1>/NM0	I0<1>/I0<1>/I0<1>/Q#6	WL<21>#1	BL#43	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<1>/NM2	I0<1>/I0<1>/I0<1>/Q#6	I0<1>/I0<1>/I0<1>/QB#3	VSS#46
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<1>/NM1	BLB#43	WL<21>#3	I0<1>/I0<1>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<1>/NM3	I0<1>/I0<1>/I0<1>/QB#4	I0<1>/I0<1>/I0<1>/Q	VSS#115
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<2>/NM0	I0<1>/I0<1>/I0<2>/Q#6	WL<22>#1	BL#41	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<2>/NM2	I0<1>/I0<1>/I0<2>/Q#6	I0<1>/I0<1>/I0<2>/QB#2	VSS#46
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<2>/NM1	BLB#43	WL<22>#4	I0<1>/I0<1>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<2>/NM3	I0<1>/I0<1>/I0<2>/QB#4	I0<1>/I0<1>/I0<2>/Q	VSS#113
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<0>/NM0	I0<1>/I0<1>/I0<0>/Q#6	WL<20>#1	BL#43	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<0>/NM2	I0<1>/I0<1>/I0<0>/Q#6	I0<1>/I0<1>/I0<0>/QB#2	VSS#48
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<1>/I0<0>/NM1	BLB#45	WL<20>#4	I0<1>/I0<1>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<1>/I0<0>/NM3	I0<1>/I0<1>/I0<0>/QB#4	I0<1>/I0<1>/I0<0>/Q	VSS#115
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<3>/NM0	I0<1>/I0<0>/I0<3>/Q#6	WL<19>#1	BL#45	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<3>/NM2	I0<1>/I0<0>/I0<3>/Q#6	I0<1>/I0<0>/I0<3>/QB#3	VSS#48
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<3>/NM1	BLB#45	WL<19>#3	I0<1>/I0<0>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<3>/NM3	I0<1>/I0<0>/I0<3>/QB#4	I0<1>/I0<0>/I0<3>/Q	VSS#117
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<1>/NM0	I0<1>/I0<0>/I0<1>/Q#6	WL<17>#1	BL#47	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<1>/NM2	I0<1>/I0<0>/I0<1>/Q#6	I0<1>/I0<0>/I0<1>/QB#3	VSS#50
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<1>/NM1	BLB#47	WL<17>#3	I0<1>/I0<0>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<1>/NM3	I0<1>/I0<0>/I0<1>/QB#4	I0<1>/I0<0>/I0<1>/Q	VSS#119
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<2>/NM0	I0<1>/I0<0>/I0<2>/Q#6	WL<18>#1	BL#45	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<2>/NM2	I0<1>/I0<0>/I0<2>/Q#6	I0<1>/I0<0>/I0<2>/QB#2	VSS#50
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<2>/NM1	BLB#47	WL<18>#4	I0<1>/I0<0>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<2>/NM3	I0<1>/I0<0>/I0<2>/QB#4	I0<1>/I0<0>/I0<2>/Q	VSS#117
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<0>/NM0	I0<1>/I0<0>/I0<0>/Q#6	WL<16>#1	BL#47	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<0>/NM2	I0<1>/I0<0>/I0<0>/Q#6	I0<1>/I0<0>/I0<0>/QB#2	VSS#52
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<1>/I0<0>/I0<0>/NM1	BLB#49	WL<16>#4	I0<1>/I0<0>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<1>/I0<0>/I0<0>/NM3	I0<1>/I0<0>/I0<0>/QB#4	I0<1>/I0<0>/I0<0>/Q	VSS#119
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<3>/NM0	I0<0>/I0<3>/I0<3>/Q#6	WL<15>#1	BL#49	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<3>/NM2	I0<0>/I0<3>/I0<3>/Q#6	I0<0>/I0<3>/I0<3>/QB#3	VSS#52
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<3>/NM1	BLB#49	WL<15>#3	I0<0>/I0<3>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<3>/NM3	I0<0>/I0<3>/I0<3>/QB#4	I0<0>/I0<3>/I0<3>/Q	VSS#121
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<1>/NM0	I0<0>/I0<3>/I0<1>/Q#6	WL<13>#1	BL#51	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<1>/NM2	I0<0>/I0<3>/I0<1>/Q#6	I0<0>/I0<3>/I0<1>/QB#3	VSS#54
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<1>/NM1	BLB#51	WL<13>#3	I0<0>/I0<3>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<1>/NM3	I0<0>/I0<3>/I0<1>/QB#4	I0<0>/I0<3>/I0<1>/Q	VSS#123
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<2>/NM0	I0<0>/I0<3>/I0<2>/Q#6	WL<14>#1	BL#49	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<2>/NM2	I0<0>/I0<3>/I0<2>/Q#6	I0<0>/I0<3>/I0<2>/QB#2	VSS#54
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<2>/NM1	BLB#51	WL<14>#4	I0<0>/I0<3>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<2>/NM3	I0<0>/I0<3>/I0<2>/QB#4	I0<0>/I0<3>/I0<2>/Q	VSS#121
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<0>/NM0	I0<0>/I0<3>/I0<0>/Q#6	WL<12>#1	BL#51	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<0>/NM2	I0<0>/I0<3>/I0<0>/Q#6	I0<0>/I0<3>/I0<0>/QB#2	VSS#56
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<3>/I0<0>/NM1	BLB#53	WL<12>#4	I0<0>/I0<3>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<3>/I0<0>/NM3	I0<0>/I0<3>/I0<0>/QB#4	I0<0>/I0<3>/I0<0>/Q	VSS#123
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<3>/NM0	I0<0>/I0<2>/I0<3>/Q#6	WL<11>#1	BL#53	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<3>/NM2	I0<0>/I0<2>/I0<3>/Q#6	I0<0>/I0<2>/I0<3>/QB#3	VSS#56
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<3>/NM1	BLB#53	WL<11>#3	I0<0>/I0<2>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<3>/NM3	I0<0>/I0<2>/I0<3>/QB#4	I0<0>/I0<2>/I0<3>/Q	VSS#125
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<1>/NM0	I0<0>/I0<2>/I0<1>/Q#6	WL<9>#1	BL#55	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<1>/NM2	I0<0>/I0<2>/I0<1>/Q#6	I0<0>/I0<2>/I0<1>/QB#3	VSS#58
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<1>/NM1	BLB#55	WL<9>#3	I0<0>/I0<2>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<1>/NM3	I0<0>/I0<2>/I0<1>/QB#4	I0<0>/I0<2>/I0<1>/Q	VSS#127
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<2>/NM0	I0<0>/I0<2>/I0<2>/Q#6	WL<10>#1	BL#53	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<2>/NM2	I0<0>/I0<2>/I0<2>/Q#6	I0<0>/I0<2>/I0<2>/QB#2	VSS#58
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<2>/NM1	BLB#55	WL<10>#4	I0<0>/I0<2>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<2>/NM3	I0<0>/I0<2>/I0<2>/QB#4	I0<0>/I0<2>/I0<2>/Q	VSS#125
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<0>/NM0	I0<0>/I0<2>/I0<0>/Q#6	WL<8>#1	BL#55	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<0>/NM2	I0<0>/I0<2>/I0<0>/Q#6	I0<0>/I0<2>/I0<0>/QB#2	VSS#60
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<2>/I0<0>/NM1	BLB#57	WL<8>#4	I0<0>/I0<2>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<2>/I0<0>/NM3	I0<0>/I0<2>/I0<0>/QB#4	I0<0>/I0<2>/I0<0>/Q	VSS#127
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<3>/NM0	I0<0>/I0<1>/I0<3>/Q#6	WL<7>#1	BL#57	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<3>/NM2	I0<0>/I0<1>/I0<3>/Q#6	I0<0>/I0<1>/I0<3>/QB#3	VSS#60
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<3>/NM1	BLB#57	WL<7>#3	I0<0>/I0<1>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<3>/NM3	I0<0>/I0<1>/I0<3>/QB#4	I0<0>/I0<1>/I0<3>/Q	VSS#129
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<1>/NM0	I0<0>/I0<1>/I0<1>/Q#6	WL<5>#1	BL#59	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<1>/NM2	I0<0>/I0<1>/I0<1>/Q#6	I0<0>/I0<1>/I0<1>/QB#3	VSS#62
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<1>/NM1	BLB#59	WL<5>#3	I0<0>/I0<1>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<1>/NM3	I0<0>/I0<1>/I0<1>/QB#4	I0<0>/I0<1>/I0<1>/Q	VSS#131
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<2>/NM0	I0<0>/I0<1>/I0<2>/Q#6	WL<6>#1	BL#57	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<2>/NM2	I0<0>/I0<1>/I0<2>/Q#6	I0<0>/I0<1>/I0<2>/QB#2	VSS#62
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<2>/NM1	BLB#59	WL<6>#4	I0<0>/I0<1>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<2>/NM3	I0<0>/I0<1>/I0<2>/QB#4	I0<0>/I0<1>/I0<2>/Q	VSS#129
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<0>/NM0	I0<0>/I0<1>/I0<0>/Q#6	WL<4>#1	BL#59	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<0>/NM2	I0<0>/I0<1>/I0<0>/Q#6	I0<0>/I0<1>/I0<0>/QB#2	VSS#64
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<1>/I0<0>/NM1	BLB#61	WL<4>#4	I0<0>/I0<1>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<1>/I0<0>/NM3	I0<0>/I0<1>/I0<0>/QB#4	I0<0>/I0<1>/I0<0>/Q	VSS#131
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<3>/NM0	I0<0>/I0<0>/I0<3>/Q#6	WL<3>#1	BL#61	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<3>/NM2	I0<0>/I0<0>/I0<3>/Q#6	I0<0>/I0<0>/I0<3>/QB#3	VSS#64
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<3>/NM1	BLB#61	WL<3>#3	I0<0>/I0<0>/I0<3>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<3>/NM3	I0<0>/I0<0>/I0<3>/QB#4	I0<0>/I0<0>/I0<3>/Q	VSS#133
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<1>/NM0	I0<0>/I0<0>/I0<1>/Q#6	WL<1>#1	BL#63	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<1>/NM2	I0<0>/I0<0>/I0<1>/Q#6	I0<0>/I0<0>/I0<1>/QB#3	VSS#66
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<1>/NM1	BLB#63	WL<1>#3	I0<0>/I0<0>/I0<1>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<1>/NM3	I0<0>/I0<0>/I0<1>/QB#4	I0<0>/I0<0>/I0<1>/Q	VSS#135
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<2>/NM0	I0<0>/I0<0>/I0<2>/Q#6	WL<2>#1	BL#61	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<2>/NM2	I0<0>/I0<0>/I0<2>/Q#6	I0<0>/I0<0>/I0<2>/QB#2	VSS#66
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<2>/NM1	BLB#63	WL<2>#4	I0<0>/I0<0>/I0<2>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<2>/NM3	I0<0>/I0<0>/I0<2>/QB#4	I0<0>/I0<0>/I0<2>/Q	VSS#133
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<0>/I0<0>/I0<0>/NM0	I0<0>/I0<0>/I0<0>/Q#6	WL<0>#1	BL#63	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.87e-14	AS=2.87e-14	PD=7e-07	PS=7e-07
MI0<0>/I0<0>/I0<0>/NM2	I0<0>/I0<0>/I0<0>/Q#6	I0<0>/I0<0>/I0<0>/QB#2	VSS#68
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I0<0>/I0<0>/NM1	BLB#65	WL<0>#4	I0<0>/I0<0>/I0<0>/QB#4	VSS#1
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I0<0>/I0<0>/NM3	I0<0>/I0<0>/I0<0>/QB#4	I0<0>/I0<0>/I0<0>/Q	VSS#135
+ VSS#1	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.75e-14	AS=3.75e-14	PD=8.1e-07	PS=8.1e-07
MI0<3>/I0<3>/I0<3>/PM0	I0<3>/I0<3>/I0<3>/Q#4	I0<3>/I0<3>/I0<3>/QB#2	VDD#2
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I0<3>/I0<3>/PM1	I0<3>/I0<3>/I0<3>/QB#5	I0<3>/I0<3>/I0<3>/Q#2	VDD#70
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<1>/PM0	I0<3>/I0<3>/I0<1>/Q#4	I0<3>/I0<3>/I0<1>/QB#2	VDD#4
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<1>/PM1	I0<3>/I0<3>/I0<1>/QB#5	I0<3>/I0<3>/I0<1>/Q#2	VDD#72
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<2>/PM0	I0<3>/I0<3>/I0<2>/Q#4	I0<3>/I0<3>/I0<2>/QB	VDD#4
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<2>/PM1	I0<3>/I0<3>/I0<2>/QB#5	I0<3>/I0<3>/I0<2>/Q#2	VDD#70
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<0>/PM0	I0<3>/I0<3>/I0<0>/Q#4	I0<3>/I0<3>/I0<0>/QB	VDD#6
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<3>/I0<0>/PM1	I0<3>/I0<3>/I0<0>/QB#5	I0<3>/I0<3>/I0<0>/Q#2	VDD#72
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<3>/PM0	I0<3>/I0<2>/I0<3>/Q#4	I0<3>/I0<2>/I0<3>/QB#2	VDD#6
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<3>/PM1	I0<3>/I0<2>/I0<3>/QB#5	I0<3>/I0<2>/I0<3>/Q#2	VDD#74
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<1>/PM0	I0<3>/I0<2>/I0<1>/Q#4	I0<3>/I0<2>/I0<1>/QB#2	VDD#8
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<1>/PM1	I0<3>/I0<2>/I0<1>/QB#5	I0<3>/I0<2>/I0<1>/Q#2	VDD#76
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<2>/PM0	I0<3>/I0<2>/I0<2>/Q#4	I0<3>/I0<2>/I0<2>/QB	VDD#8
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<2>/PM1	I0<3>/I0<2>/I0<2>/QB#5	I0<3>/I0<2>/I0<2>/Q#2	VDD#74
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<0>/PM0	I0<3>/I0<2>/I0<0>/Q#4	I0<3>/I0<2>/I0<0>/QB	VDD#10
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<2>/I0<0>/PM1	I0<3>/I0<2>/I0<0>/QB#5	I0<3>/I0<2>/I0<0>/Q#2	VDD#76
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<3>/PM0	I0<3>/I0<1>/I0<3>/Q#4	I0<3>/I0<1>/I0<3>/QB#2	VDD#10
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<3>/PM1	I0<3>/I0<1>/I0<3>/QB#5	I0<3>/I0<1>/I0<3>/Q#2	VDD#78
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<1>/PM0	I0<3>/I0<1>/I0<1>/Q#4	I0<3>/I0<1>/I0<1>/QB#2	VDD#12
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<1>/PM1	I0<3>/I0<1>/I0<1>/QB#5	I0<3>/I0<1>/I0<1>/Q#2	VDD#80
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<2>/PM0	I0<3>/I0<1>/I0<2>/Q#4	I0<3>/I0<1>/I0<2>/QB	VDD#12
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<2>/PM1	I0<3>/I0<1>/I0<2>/QB#5	I0<3>/I0<1>/I0<2>/Q#2	VDD#78
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<0>/PM0	I0<3>/I0<1>/I0<0>/Q#4	I0<3>/I0<1>/I0<0>/QB	VDD#14
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<1>/I0<0>/PM1	I0<3>/I0<1>/I0<0>/QB#5	I0<3>/I0<1>/I0<0>/Q#2	VDD#80
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<3>/PM0	I0<3>/I0<0>/I0<3>/Q#4	I0<3>/I0<0>/I0<3>/QB#2	VDD#14
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<3>/PM1	I0<3>/I0<0>/I0<3>/QB#5	I0<3>/I0<0>/I0<3>/Q#2	VDD#82
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<1>/PM0	I0<3>/I0<0>/I0<1>/Q#4	I0<3>/I0<0>/I0<1>/QB#2	VDD#16
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<1>/PM1	I0<3>/I0<0>/I0<1>/QB#5	I0<3>/I0<0>/I0<1>/Q#2	VDD#84
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<2>/PM0	I0<3>/I0<0>/I0<2>/Q#4	I0<3>/I0<0>/I0<2>/QB	VDD#16
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<2>/PM1	I0<3>/I0<0>/I0<2>/QB#5	I0<3>/I0<0>/I0<2>/Q#2	VDD#82
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<0>/PM0	I0<3>/I0<0>/I0<0>/Q#4	I0<3>/I0<0>/I0<0>/QB	VDD#18
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<3>/I0<0>/I0<0>/PM1	I0<3>/I0<0>/I0<0>/QB#5	I0<3>/I0<0>/I0<0>/Q#2	VDD#84
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<3>/PM0	I0<2>/I0<3>/I0<3>/Q#4	I0<2>/I0<3>/I0<3>/QB#2	VDD#18
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<3>/PM1	I0<2>/I0<3>/I0<3>/QB#5	I0<2>/I0<3>/I0<3>/Q#2	VDD#86
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<1>/PM0	I0<2>/I0<3>/I0<1>/Q#4	I0<2>/I0<3>/I0<1>/QB#2	VDD#20
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<1>/PM1	I0<2>/I0<3>/I0<1>/QB#5	I0<2>/I0<3>/I0<1>/Q#2	VDD#88
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<2>/PM0	I0<2>/I0<3>/I0<2>/Q#4	I0<2>/I0<3>/I0<2>/QB	VDD#20
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<2>/PM1	I0<2>/I0<3>/I0<2>/QB#5	I0<2>/I0<3>/I0<2>/Q#2	VDD#86
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<0>/PM0	I0<2>/I0<3>/I0<0>/Q#4	I0<2>/I0<3>/I0<0>/QB	VDD#22
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<3>/I0<0>/PM1	I0<2>/I0<3>/I0<0>/QB#5	I0<2>/I0<3>/I0<0>/Q#2	VDD#88
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<3>/PM0	I0<2>/I0<2>/I0<3>/Q#4	I0<2>/I0<2>/I0<3>/QB#2	VDD#22
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<3>/PM1	I0<2>/I0<2>/I0<3>/QB#5	I0<2>/I0<2>/I0<3>/Q#2	VDD#90
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<1>/PM0	I0<2>/I0<2>/I0<1>/Q#4	I0<2>/I0<2>/I0<1>/QB#2	VDD#24
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<1>/PM1	I0<2>/I0<2>/I0<1>/QB#5	I0<2>/I0<2>/I0<1>/Q#2	VDD#92
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<2>/PM0	I0<2>/I0<2>/I0<2>/Q#4	I0<2>/I0<2>/I0<2>/QB	VDD#24
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<2>/PM1	I0<2>/I0<2>/I0<2>/QB#5	I0<2>/I0<2>/I0<2>/Q#2	VDD#90
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<0>/PM0	I0<2>/I0<2>/I0<0>/Q#4	I0<2>/I0<2>/I0<0>/QB	VDD#26
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<2>/I0<0>/PM1	I0<2>/I0<2>/I0<0>/QB#5	I0<2>/I0<2>/I0<0>/Q#2	VDD#92
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<3>/PM0	I0<2>/I0<1>/I0<3>/Q#4	I0<2>/I0<1>/I0<3>/QB#2	VDD#26
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<3>/PM1	I0<2>/I0<1>/I0<3>/QB#5	I0<2>/I0<1>/I0<3>/Q#2	VDD#94
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<1>/PM0	I0<2>/I0<1>/I0<1>/Q#4	I0<2>/I0<1>/I0<1>/QB#2	VDD#28
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<1>/PM1	I0<2>/I0<1>/I0<1>/QB#5	I0<2>/I0<1>/I0<1>/Q#2	VDD#96
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<2>/PM0	I0<2>/I0<1>/I0<2>/Q#4	I0<2>/I0<1>/I0<2>/QB	VDD#28
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<2>/PM1	I0<2>/I0<1>/I0<2>/QB#5	I0<2>/I0<1>/I0<2>/Q#2	VDD#94
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<0>/PM0	I0<2>/I0<1>/I0<0>/Q#4	I0<2>/I0<1>/I0<0>/QB	VDD#30
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<1>/I0<0>/PM1	I0<2>/I0<1>/I0<0>/QB#5	I0<2>/I0<1>/I0<0>/Q#2	VDD#96
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<3>/PM0	I0<2>/I0<0>/I0<3>/Q#4	I0<2>/I0<0>/I0<3>/QB#2	VDD#30
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<3>/PM1	I0<2>/I0<0>/I0<3>/QB#5	I0<2>/I0<0>/I0<3>/Q#2	VDD#98
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<1>/PM0	I0<2>/I0<0>/I0<1>/Q#4	I0<2>/I0<0>/I0<1>/QB#2	VDD#32
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<1>/PM1	I0<2>/I0<0>/I0<1>/QB#5	I0<2>/I0<0>/I0<1>/Q#2	VDD#100
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<2>/PM0	I0<2>/I0<0>/I0<2>/Q#4	I0<2>/I0<0>/I0<2>/QB	VDD#32
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<2>/PM1	I0<2>/I0<0>/I0<2>/QB#5	I0<2>/I0<0>/I0<2>/Q#2	VDD#98
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<0>/PM0	I0<2>/I0<0>/I0<0>/Q#4	I0<2>/I0<0>/I0<0>/QB	VDD#34
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<2>/I0<0>/I0<0>/PM1	I0<2>/I0<0>/I0<0>/QB#5	I0<2>/I0<0>/I0<0>/Q#2	VDD#100
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<3>/PM0	I0<1>/I0<3>/I0<3>/Q#4	I0<1>/I0<3>/I0<3>/QB#2	VDD#34
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<3>/PM1	I0<1>/I0<3>/I0<3>/QB#5	I0<1>/I0<3>/I0<3>/Q#2	VDD#102
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<1>/PM0	I0<1>/I0<3>/I0<1>/Q#4	I0<1>/I0<3>/I0<1>/QB#2	VDD#36
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<1>/PM1	I0<1>/I0<3>/I0<1>/QB#5	I0<1>/I0<3>/I0<1>/Q#2	VDD#104
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<2>/PM0	I0<1>/I0<3>/I0<2>/Q#4	I0<1>/I0<3>/I0<2>/QB	VDD#36
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<2>/PM1	I0<1>/I0<3>/I0<2>/QB#5	I0<1>/I0<3>/I0<2>/Q#2	VDD#102
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<0>/PM0	I0<1>/I0<3>/I0<0>/Q#4	I0<1>/I0<3>/I0<0>/QB	VDD#38
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<3>/I0<0>/PM1	I0<1>/I0<3>/I0<0>/QB#5	I0<1>/I0<3>/I0<0>/Q#2	VDD#104
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<3>/PM0	I0<1>/I0<2>/I0<3>/Q#4	I0<1>/I0<2>/I0<3>/QB#2	VDD#38
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<3>/PM1	I0<1>/I0<2>/I0<3>/QB#5	I0<1>/I0<2>/I0<3>/Q#2	VDD#106
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<1>/PM0	I0<1>/I0<2>/I0<1>/Q#4	I0<1>/I0<2>/I0<1>/QB#2	VDD#40
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<1>/PM1	I0<1>/I0<2>/I0<1>/QB#5	I0<1>/I0<2>/I0<1>/Q#2	VDD#108
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<2>/PM0	I0<1>/I0<2>/I0<2>/Q#4	I0<1>/I0<2>/I0<2>/QB	VDD#40
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<2>/PM1	I0<1>/I0<2>/I0<2>/QB#5	I0<1>/I0<2>/I0<2>/Q#2	VDD#106
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<0>/PM0	I0<1>/I0<2>/I0<0>/Q#4	I0<1>/I0<2>/I0<0>/QB	VDD#42
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<2>/I0<0>/PM1	I0<1>/I0<2>/I0<0>/QB#5	I0<1>/I0<2>/I0<0>/Q#2	VDD#108
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<3>/PM0	I0<1>/I0<1>/I0<3>/Q#4	I0<1>/I0<1>/I0<3>/QB#2	VDD#42
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<3>/PM1	I0<1>/I0<1>/I0<3>/QB#5	I0<1>/I0<1>/I0<3>/Q#2	VDD#110
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<1>/PM0	I0<1>/I0<1>/I0<1>/Q#4	I0<1>/I0<1>/I0<1>/QB#2	VDD#44
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<1>/PM1	I0<1>/I0<1>/I0<1>/QB#5	I0<1>/I0<1>/I0<1>/Q#2	VDD#112
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<2>/PM0	I0<1>/I0<1>/I0<2>/Q#4	I0<1>/I0<1>/I0<2>/QB	VDD#44
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<2>/PM1	I0<1>/I0<1>/I0<2>/QB#5	I0<1>/I0<1>/I0<2>/Q#2	VDD#110
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<0>/PM0	I0<1>/I0<1>/I0<0>/Q#4	I0<1>/I0<1>/I0<0>/QB	VDD#46
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<1>/I0<0>/PM1	I0<1>/I0<1>/I0<0>/QB#5	I0<1>/I0<1>/I0<0>/Q#2	VDD#112
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<3>/PM0	I0<1>/I0<0>/I0<3>/Q#4	I0<1>/I0<0>/I0<3>/QB#2	VDD#46
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<3>/PM1	I0<1>/I0<0>/I0<3>/QB#5	I0<1>/I0<0>/I0<3>/Q#2	VDD#114
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<1>/PM0	I0<1>/I0<0>/I0<1>/Q#4	I0<1>/I0<0>/I0<1>/QB#2	VDD#48
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<1>/PM1	I0<1>/I0<0>/I0<1>/QB#5	I0<1>/I0<0>/I0<1>/Q#2	VDD#116
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<2>/PM0	I0<1>/I0<0>/I0<2>/Q#4	I0<1>/I0<0>/I0<2>/QB	VDD#48
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<2>/PM1	I0<1>/I0<0>/I0<2>/QB#5	I0<1>/I0<0>/I0<2>/Q#2	VDD#114
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<0>/PM0	I0<1>/I0<0>/I0<0>/Q#4	I0<1>/I0<0>/I0<0>/QB	VDD#50
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<1>/I0<0>/I0<0>/PM1	I0<1>/I0<0>/I0<0>/QB#5	I0<1>/I0<0>/I0<0>/Q#2	VDD#116
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<3>/PM0	I0<0>/I0<3>/I0<3>/Q#4	I0<0>/I0<3>/I0<3>/QB#2	VDD#50
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<3>/PM1	I0<0>/I0<3>/I0<3>/QB#5	I0<0>/I0<3>/I0<3>/Q#2	VDD#118
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<1>/PM0	I0<0>/I0<3>/I0<1>/Q#4	I0<0>/I0<3>/I0<1>/QB#2	VDD#52
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<1>/PM1	I0<0>/I0<3>/I0<1>/QB#5	I0<0>/I0<3>/I0<1>/Q#2	VDD#120
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<2>/PM0	I0<0>/I0<3>/I0<2>/Q#4	I0<0>/I0<3>/I0<2>/QB	VDD#52
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<2>/PM1	I0<0>/I0<3>/I0<2>/QB#5	I0<0>/I0<3>/I0<2>/Q#2	VDD#118
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<0>/PM0	I0<0>/I0<3>/I0<0>/Q#4	I0<0>/I0<3>/I0<0>/QB	VDD#54
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<3>/I0<0>/PM1	I0<0>/I0<3>/I0<0>/QB#5	I0<0>/I0<3>/I0<0>/Q#2	VDD#120
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<3>/PM0	I0<0>/I0<2>/I0<3>/Q#4	I0<0>/I0<2>/I0<3>/QB#2	VDD#54
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<3>/PM1	I0<0>/I0<2>/I0<3>/QB#5	I0<0>/I0<2>/I0<3>/Q#2	VDD#122
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<1>/PM0	I0<0>/I0<2>/I0<1>/Q#4	I0<0>/I0<2>/I0<1>/QB#2	VDD#56
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<1>/PM1	I0<0>/I0<2>/I0<1>/QB#5	I0<0>/I0<2>/I0<1>/Q#2	VDD#124
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<2>/PM0	I0<0>/I0<2>/I0<2>/Q#4	I0<0>/I0<2>/I0<2>/QB	VDD#56
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<2>/PM1	I0<0>/I0<2>/I0<2>/QB#5	I0<0>/I0<2>/I0<2>/Q#2	VDD#122
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<0>/PM0	I0<0>/I0<2>/I0<0>/Q#4	I0<0>/I0<2>/I0<0>/QB	VDD#58
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<2>/I0<0>/PM1	I0<0>/I0<2>/I0<0>/QB#5	I0<0>/I0<2>/I0<0>/Q#2	VDD#124
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<3>/PM0	I0<0>/I0<1>/I0<3>/Q#4	I0<0>/I0<1>/I0<3>/QB#2	VDD#58
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<3>/PM1	I0<0>/I0<1>/I0<3>/QB#5	I0<0>/I0<1>/I0<3>/Q#2	VDD#126
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<1>/PM0	I0<0>/I0<1>/I0<1>/Q#4	I0<0>/I0<1>/I0<1>/QB#2	VDD#60
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<1>/PM1	I0<0>/I0<1>/I0<1>/QB#5	I0<0>/I0<1>/I0<1>/Q#2	VDD#128
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<2>/PM0	I0<0>/I0<1>/I0<2>/Q#4	I0<0>/I0<1>/I0<2>/QB	VDD#60
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<2>/PM1	I0<0>/I0<1>/I0<2>/QB#5	I0<0>/I0<1>/I0<2>/Q#2	VDD#126
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<0>/PM0	I0<0>/I0<1>/I0<0>/Q#4	I0<0>/I0<1>/I0<0>/QB	VDD#62
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<1>/I0<0>/PM1	I0<0>/I0<1>/I0<0>/QB#5	I0<0>/I0<1>/I0<0>/Q#2	VDD#128
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<3>/PM0	I0<0>/I0<0>/I0<3>/Q#4	I0<0>/I0<0>/I0<3>/QB#2	VDD#62
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<3>/PM1	I0<0>/I0<0>/I0<3>/QB#5	I0<0>/I0<0>/I0<3>/Q#2	VDD#130
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<1>/PM0	I0<0>/I0<0>/I0<1>/Q#4	I0<0>/I0<0>/I0<1>/QB#2	VDD#64
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<1>/PM1	I0<0>/I0<0>/I0<1>/QB#5	I0<0>/I0<0>/I0<1>/Q#2	VDD#132
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<2>/PM0	I0<0>/I0<0>/I0<2>/Q#4	I0<0>/I0<0>/I0<2>/QB	VDD#64
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<2>/PM1	I0<0>/I0<0>/I0<2>/QB#5	I0<0>/I0<0>/I0<2>/Q#2	VDD#130
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
MI0<0>/I0<0>/I0<0>/PM0	I0<0>/I0<0>/I0<0>/Q#4	I0<0>/I0<0>/I0<0>/QB	VDD#66
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I0<0>/I0<0>/PM1	I0<0>/I0<0>/I0<0>/QB#5	I0<0>/I0<0>/I0<0>/Q#2	VDD#132
+ VDD#68	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.8e-14	AS=1.8e-14	PD=5.4e-07	PS=5.4e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	WL<63>#1	WL<63>#2	  104.7064	$poly_conn
Rl2	WL<62>#1	WL<62>#2	  104.7064	$poly_conn
Rl3	WL<61>#1	WL<61>#2	  104.7064	$poly_conn
Rl4	WL<60>#1	WL<60>#2	  104.7064	$poly_conn
Rl5	WL<59>#1	WL<59>#2	  104.7064	$poly_conn
Rl6	WL<58>#1	WL<58>#2	  104.7064	$poly_conn
Rl7	WL<57>#1	WL<57>#2	  104.7064	$poly_conn
Rl8	WL<56>#1	WL<56>#2	  104.7064	$poly_conn
Rl9	WL<55>#1	WL<55>#2	  104.7064	$poly_conn
Rl10	WL<54>#1	WL<54>#2	  104.7064	$poly_conn
Rl11	WL<53>#1	WL<53>#2	  104.7064	$poly_conn
Rl12	WL<52>#1	WL<52>#2	  104.7064	$poly_conn
Rl13	WL<51>#1	WL<51>#2	  104.7064	$poly_conn
Rl14	WL<50>#1	WL<50>#2	  104.7064	$poly_conn
Rl15	WL<49>#1	WL<49>#2	  104.7064	$poly_conn
Rl16	WL<48>#1	WL<48>#2	  104.7064	$poly_conn
Rl17	WL<47>#1	WL<47>#2	  104.7064	$poly_conn
Rl18	WL<46>#1	WL<46>#2	  104.7064	$poly_conn
Rl19	WL<45>#1	WL<45>#2	  104.7064	$poly_conn
Rl20	WL<44>#1	WL<44>#2	  104.7064	$poly_conn
Rl21	WL<43>#1	WL<43>#2	  104.7064	$poly_conn
Rl22	WL<42>#1	WL<42>#2	  104.7064	$poly_conn
Rl23	WL<41>#1	WL<41>#2	  104.7064	$poly_conn
Rl24	WL<40>#1	WL<40>#2	  104.7064	$poly_conn
Rl25	WL<39>#1	WL<39>#2	  104.7064	$poly_conn
Rl26	WL<38>#1	WL<38>#2	  104.7064	$poly_conn
Rl27	WL<37>#1	WL<37>#2	  104.7064	$poly_conn
Rl28	WL<36>#1	WL<36>#2	  104.7064	$poly_conn
Rl29	WL<35>#1	WL<35>#2	  104.7064	$poly_conn
Rl30	WL<34>#1	WL<34>#2	  104.7064	$poly_conn
Rl31	WL<33>#1	WL<33>#2	  104.7064	$poly_conn
Rl32	WL<32>#1	WL<32>#2	  104.7064	$poly_conn
Rl33	WL<31>#1	WL<31>#2	  104.7064	$poly_conn
Rl34	WL<30>#1	WL<30>#2	  104.7064	$poly_conn
Rl35	WL<29>#1	WL<29>#2	  104.7064	$poly_conn
Rl36	WL<28>#1	WL<28>#2	  104.7064	$poly_conn
Rl37	WL<27>#1	WL<27>#2	  104.7064	$poly_conn
Rl38	WL<26>#1	WL<26>#2	  104.7064	$poly_conn
Rl39	WL<25>#1	WL<25>#2	  104.7064	$poly_conn
Rl40	WL<24>#1	WL<24>#2	  104.7064	$poly_conn
Rl41	WL<23>#1	WL<23>#2	  104.7064	$poly_conn
Rl42	WL<22>#1	WL<22>#2	  104.7064	$poly_conn
Rl43	WL<21>#1	WL<21>#2	  104.7064	$poly_conn
Rl44	WL<20>#1	WL<20>#2	  104.7064	$poly_conn
Rl45	WL<19>#1	WL<19>#2	  104.7064	$poly_conn
Rl46	WL<18>#1	WL<18>#2	  104.7064	$poly_conn
Rl47	WL<17>#1	WL<17>#2	  104.7064	$poly_conn
Rl48	WL<16>#1	WL<16>#2	  104.7064	$poly_conn
Rl49	WL<15>#1	WL<15>#2	  104.7064	$poly_conn
Rl50	WL<14>#1	WL<14>#2	  104.7064	$poly_conn
Rl51	WL<13>#1	WL<13>#2	  104.7064	$poly_conn
Rl52	WL<12>#1	WL<12>#2	  104.7064	$poly_conn
Rl53	WL<11>#1	WL<11>#2	  104.7064	$poly_conn
Rl54	WL<10>#1	WL<10>#2	  104.7064	$poly_conn
Rl55	WL<9>#1	WL<9>#2	  104.7064	$poly_conn
Rl56	WL<8>#1	WL<8>#2	  104.7064	$poly_conn
Rl57	WL<7>#1	WL<7>#2	  104.7064	$poly_conn
Rl58	WL<6>#1	WL<6>#2	  104.7064	$poly_conn
Rl59	WL<5>#1	WL<5>#2	  104.7064	$poly_conn
Rl60	WL<4>#1	WL<4>#2	  104.7064	$poly_conn
Rl61	WL<3>#1	WL<3>#2	  104.7064	$poly_conn
Rl62	WL<2>#1	WL<2>#2	  104.7064	$poly_conn
Rl63	WL<1>#1	WL<1>#2	  104.7064	$poly_conn
Rl64	WL<0>#1	WL<0>#2	  104.7064	$poly_conn
Rl65	I0<3>/I0<3>/I0<3>/QB	I0<3>/I0<3>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl66	I0<3>/I0<3>/I0<3>/QB#2	I0<3>/I0<3>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl67	I0<3>/I0<3>/I0<2>/QB	I0<3>/I0<3>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl68	I0<3>/I0<3>/I0<2>/QB	I0<3>/I0<3>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl69	I0<3>/I0<3>/I0<1>/QB	I0<3>/I0<3>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl70	I0<3>/I0<3>/I0<1>/QB#2	I0<3>/I0<3>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl71	I0<3>/I0<3>/I0<0>/QB	I0<3>/I0<3>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl72	I0<3>/I0<3>/I0<0>/QB	I0<3>/I0<3>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl73	I0<3>/I0<2>/I0<3>/QB	I0<3>/I0<2>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl74	I0<3>/I0<2>/I0<3>/QB#2	I0<3>/I0<2>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl75	I0<3>/I0<2>/I0<2>/QB	I0<3>/I0<2>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl76	I0<3>/I0<2>/I0<2>/QB	I0<3>/I0<2>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl77	I0<3>/I0<2>/I0<1>/QB	I0<3>/I0<2>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl78	I0<3>/I0<2>/I0<1>/QB#2	I0<3>/I0<2>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl79	I0<3>/I0<2>/I0<0>/QB	I0<3>/I0<2>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl80	I0<3>/I0<2>/I0<0>/QB	I0<3>/I0<2>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl81	I0<3>/I0<1>/I0<3>/QB	I0<3>/I0<1>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl82	I0<3>/I0<1>/I0<3>/QB#2	I0<3>/I0<1>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl83	I0<3>/I0<1>/I0<2>/QB	I0<3>/I0<1>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl84	I0<3>/I0<1>/I0<2>/QB	I0<3>/I0<1>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl85	I0<3>/I0<1>/I0<1>/QB	I0<3>/I0<1>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl86	I0<3>/I0<1>/I0<1>/QB#2	I0<3>/I0<1>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl87	I0<3>/I0<1>/I0<0>/QB	I0<3>/I0<1>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl88	I0<3>/I0<1>/I0<0>/QB	I0<3>/I0<1>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl89	I0<3>/I0<0>/I0<3>/QB	I0<3>/I0<0>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl90	I0<3>/I0<0>/I0<3>/QB#2	I0<3>/I0<0>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl91	I0<3>/I0<0>/I0<2>/QB	I0<3>/I0<0>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl92	I0<3>/I0<0>/I0<2>/QB	I0<3>/I0<0>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl93	I0<3>/I0<0>/I0<1>/QB	I0<3>/I0<0>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl94	I0<3>/I0<0>/I0<1>/QB#2	I0<3>/I0<0>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl95	I0<3>/I0<0>/I0<0>/QB	I0<3>/I0<0>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl96	I0<3>/I0<0>/I0<0>/QB	I0<3>/I0<0>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl97	I0<2>/I0<3>/I0<3>/QB	I0<2>/I0<3>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl98	I0<2>/I0<3>/I0<3>/QB#2	I0<2>/I0<3>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl99	I0<2>/I0<3>/I0<2>/QB	I0<2>/I0<3>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl100	I0<2>/I0<3>/I0<2>/QB	I0<2>/I0<3>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl101	I0<2>/I0<3>/I0<1>/QB	I0<2>/I0<3>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl102	I0<2>/I0<3>/I0<1>/QB#2	I0<2>/I0<3>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl103	I0<2>/I0<3>/I0<0>/QB	I0<2>/I0<3>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl104	I0<2>/I0<3>/I0<0>/QB	I0<2>/I0<3>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl105	I0<2>/I0<2>/I0<3>/QB	I0<2>/I0<2>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl106	I0<2>/I0<2>/I0<3>/QB#2	I0<2>/I0<2>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl107	I0<2>/I0<2>/I0<2>/QB	I0<2>/I0<2>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl108	I0<2>/I0<2>/I0<2>/QB	I0<2>/I0<2>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl109	I0<2>/I0<2>/I0<1>/QB	I0<2>/I0<2>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl110	I0<2>/I0<2>/I0<1>/QB#2	I0<2>/I0<2>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl111	I0<2>/I0<2>/I0<0>/QB	I0<2>/I0<2>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl112	I0<2>/I0<2>/I0<0>/QB	I0<2>/I0<2>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl113	I0<2>/I0<1>/I0<3>/QB	I0<2>/I0<1>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl114	I0<2>/I0<1>/I0<3>/QB#2	I0<2>/I0<1>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl115	I0<2>/I0<1>/I0<2>/QB	I0<2>/I0<1>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl116	I0<2>/I0<1>/I0<2>/QB	I0<2>/I0<1>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl117	I0<2>/I0<1>/I0<1>/QB	I0<2>/I0<1>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl118	I0<2>/I0<1>/I0<1>/QB#2	I0<2>/I0<1>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl119	I0<2>/I0<1>/I0<0>/QB	I0<2>/I0<1>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl120	I0<2>/I0<1>/I0<0>/QB	I0<2>/I0<1>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl121	I0<2>/I0<0>/I0<3>/QB	I0<2>/I0<0>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl122	I0<2>/I0<0>/I0<3>/QB#2	I0<2>/I0<0>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl123	I0<2>/I0<0>/I0<2>/QB	I0<2>/I0<0>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl124	I0<2>/I0<0>/I0<2>/QB	I0<2>/I0<0>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl125	I0<2>/I0<0>/I0<1>/QB	I0<2>/I0<0>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl126	I0<2>/I0<0>/I0<1>/QB#2	I0<2>/I0<0>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl127	I0<2>/I0<0>/I0<0>/QB	I0<2>/I0<0>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl128	I0<2>/I0<0>/I0<0>/QB	I0<2>/I0<0>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl129	I0<1>/I0<3>/I0<3>/QB	I0<1>/I0<3>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl130	I0<1>/I0<3>/I0<3>/QB#2	I0<1>/I0<3>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl131	I0<1>/I0<3>/I0<2>/QB	I0<1>/I0<3>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl132	I0<1>/I0<3>/I0<2>/QB	I0<1>/I0<3>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl133	I0<1>/I0<3>/I0<1>/QB	I0<1>/I0<3>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl134	I0<1>/I0<3>/I0<1>/QB#2	I0<1>/I0<3>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl135	I0<1>/I0<3>/I0<0>/QB	I0<1>/I0<3>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl136	I0<1>/I0<3>/I0<0>/QB	I0<1>/I0<3>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl137	I0<1>/I0<2>/I0<3>/QB	I0<1>/I0<2>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl138	I0<1>/I0<2>/I0<3>/QB#2	I0<1>/I0<2>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl139	I0<1>/I0<2>/I0<2>/QB	I0<1>/I0<2>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl140	I0<1>/I0<2>/I0<2>/QB	I0<1>/I0<2>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl141	I0<1>/I0<2>/I0<1>/QB	I0<1>/I0<2>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl142	I0<1>/I0<2>/I0<1>/QB#2	I0<1>/I0<2>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl143	I0<1>/I0<2>/I0<0>/QB	I0<1>/I0<2>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl144	I0<1>/I0<2>/I0<0>/QB	I0<1>/I0<2>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl145	I0<1>/I0<1>/I0<3>/QB	I0<1>/I0<1>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl146	I0<1>/I0<1>/I0<3>/QB#2	I0<1>/I0<1>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl147	I0<1>/I0<1>/I0<2>/QB	I0<1>/I0<1>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl148	I0<1>/I0<1>/I0<2>/QB	I0<1>/I0<1>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl149	I0<1>/I0<1>/I0<1>/QB	I0<1>/I0<1>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl150	I0<1>/I0<1>/I0<1>/QB#2	I0<1>/I0<1>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl151	I0<1>/I0<1>/I0<0>/QB	I0<1>/I0<1>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl152	I0<1>/I0<1>/I0<0>/QB	I0<1>/I0<1>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl153	I0<1>/I0<0>/I0<3>/QB	I0<1>/I0<0>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl154	I0<1>/I0<0>/I0<3>/QB#2	I0<1>/I0<0>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl155	I0<1>/I0<0>/I0<2>/QB	I0<1>/I0<0>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl156	I0<1>/I0<0>/I0<2>/QB	I0<1>/I0<0>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl157	I0<1>/I0<0>/I0<1>/QB	I0<1>/I0<0>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl158	I0<1>/I0<0>/I0<1>/QB#2	I0<1>/I0<0>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl159	I0<1>/I0<0>/I0<0>/QB	I0<1>/I0<0>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl160	I0<1>/I0<0>/I0<0>/QB	I0<1>/I0<0>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl161	I0<0>/I0<3>/I0<3>/QB	I0<0>/I0<3>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl162	I0<0>/I0<3>/I0<3>/QB#2	I0<0>/I0<3>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl163	I0<0>/I0<3>/I0<2>/QB	I0<0>/I0<3>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl164	I0<0>/I0<3>/I0<2>/QB	I0<0>/I0<3>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl165	I0<0>/I0<3>/I0<1>/QB	I0<0>/I0<3>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl166	I0<0>/I0<3>/I0<1>/QB#2	I0<0>/I0<3>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl167	I0<0>/I0<3>/I0<0>/QB	I0<0>/I0<3>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl168	I0<0>/I0<3>/I0<0>/QB	I0<0>/I0<3>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl169	I0<0>/I0<2>/I0<3>/QB	I0<0>/I0<2>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl170	I0<0>/I0<2>/I0<3>/QB#2	I0<0>/I0<2>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl171	I0<0>/I0<2>/I0<2>/QB	I0<0>/I0<2>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl172	I0<0>/I0<2>/I0<2>/QB	I0<0>/I0<2>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl173	I0<0>/I0<2>/I0<1>/QB	I0<0>/I0<2>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl174	I0<0>/I0<2>/I0<1>/QB#2	I0<0>/I0<2>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl175	I0<0>/I0<2>/I0<0>/QB	I0<0>/I0<2>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl176	I0<0>/I0<2>/I0<0>/QB	I0<0>/I0<2>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl177	I0<0>/I0<1>/I0<3>/QB	I0<0>/I0<1>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl178	I0<0>/I0<1>/I0<3>/QB#2	I0<0>/I0<1>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl179	I0<0>/I0<1>/I0<2>/QB	I0<0>/I0<1>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl180	I0<0>/I0<1>/I0<2>/QB	I0<0>/I0<1>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl181	I0<0>/I0<1>/I0<1>/QB	I0<0>/I0<1>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl182	I0<0>/I0<1>/I0<1>/QB#2	I0<0>/I0<1>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl183	I0<0>/I0<1>/I0<0>/QB	I0<0>/I0<1>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl184	I0<0>/I0<1>/I0<0>/QB	I0<0>/I0<1>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl185	I0<0>/I0<0>/I0<3>/QB	I0<0>/I0<0>/I0<3>/QB#2	   90.3330
+ $poly_conn
Rl186	I0<0>/I0<0>/I0<3>/QB#2	I0<0>/I0<0>/I0<3>/QB#3	   56.4103
+ $poly_conn
Rl187	I0<0>/I0<0>/I0<2>/QB	I0<0>/I0<0>/I0<2>/QB#2	   56.4103
+ $poly_conn
Rl188	I0<0>/I0<0>/I0<2>/QB	I0<0>/I0<0>/I0<2>/QB#3	   90.3330
+ $poly_conn
Rl189	I0<0>/I0<0>/I0<1>/QB	I0<0>/I0<0>/I0<1>/QB#2	   90.3330
+ $poly_conn
Rl190	I0<0>/I0<0>/I0<1>/QB#2	I0<0>/I0<0>/I0<1>/QB#3	   56.4103
+ $poly_conn
Rl191	I0<0>/I0<0>/I0<0>/QB	I0<0>/I0<0>/I0<0>/QB#2	   56.4103
+ $poly_conn
Rl192	I0<0>/I0<0>/I0<0>/QB	I0<0>/I0<0>/I0<0>/QB#3	   90.3330
+ $poly_conn
Rl193	I0<3>/I0<3>/I0<3>/Q	I0<3>/I0<3>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl194	I0<3>/I0<3>/I0<3>/Q#2	I0<3>/I0<3>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl195	I0<3>/I0<3>/I0<2>/Q	I0<3>/I0<3>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl196	I0<3>/I0<3>/I0<2>/Q#2	I0<3>/I0<3>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl197	I0<3>/I0<3>/I0<1>/Q	I0<3>/I0<3>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl198	I0<3>/I0<3>/I0<1>/Q#2	I0<3>/I0<3>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl199	I0<3>/I0<3>/I0<0>/Q	I0<3>/I0<3>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl200	I0<3>/I0<3>/I0<0>/Q#2	I0<3>/I0<3>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl201	I0<3>/I0<2>/I0<3>/Q	I0<3>/I0<2>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl202	I0<3>/I0<2>/I0<3>/Q#2	I0<3>/I0<2>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl203	I0<3>/I0<2>/I0<2>/Q	I0<3>/I0<2>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl204	I0<3>/I0<2>/I0<2>/Q#2	I0<3>/I0<2>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl205	I0<3>/I0<2>/I0<1>/Q	I0<3>/I0<2>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl206	I0<3>/I0<2>/I0<1>/Q#2	I0<3>/I0<2>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl207	I0<3>/I0<2>/I0<0>/Q	I0<3>/I0<2>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl208	I0<3>/I0<2>/I0<0>/Q#2	I0<3>/I0<2>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl209	I0<3>/I0<1>/I0<3>/Q	I0<3>/I0<1>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl210	I0<3>/I0<1>/I0<3>/Q#2	I0<3>/I0<1>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl211	I0<3>/I0<1>/I0<2>/Q	I0<3>/I0<1>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl212	I0<3>/I0<1>/I0<2>/Q#2	I0<3>/I0<1>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl213	I0<3>/I0<1>/I0<1>/Q	I0<3>/I0<1>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl214	I0<3>/I0<1>/I0<1>/Q#2	I0<3>/I0<1>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl215	I0<3>/I0<1>/I0<0>/Q	I0<3>/I0<1>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl216	I0<3>/I0<1>/I0<0>/Q#2	I0<3>/I0<1>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl217	I0<3>/I0<0>/I0<3>/Q	I0<3>/I0<0>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl218	I0<3>/I0<0>/I0<3>/Q#2	I0<3>/I0<0>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl219	I0<3>/I0<0>/I0<2>/Q	I0<3>/I0<0>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl220	I0<3>/I0<0>/I0<2>/Q#2	I0<3>/I0<0>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl221	I0<3>/I0<0>/I0<1>/Q	I0<3>/I0<0>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl222	I0<3>/I0<0>/I0<1>/Q#2	I0<3>/I0<0>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl223	I0<3>/I0<0>/I0<0>/Q	I0<3>/I0<0>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl224	I0<3>/I0<0>/I0<0>/Q#2	I0<3>/I0<0>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl225	I0<2>/I0<3>/I0<3>/Q	I0<2>/I0<3>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl226	I0<2>/I0<3>/I0<3>/Q#2	I0<2>/I0<3>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl227	I0<2>/I0<3>/I0<2>/Q	I0<2>/I0<3>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl228	I0<2>/I0<3>/I0<2>/Q#2	I0<2>/I0<3>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl229	I0<2>/I0<3>/I0<1>/Q	I0<2>/I0<3>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl230	I0<2>/I0<3>/I0<1>/Q#2	I0<2>/I0<3>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl231	I0<2>/I0<3>/I0<0>/Q	I0<2>/I0<3>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl232	I0<2>/I0<3>/I0<0>/Q#2	I0<2>/I0<3>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl233	I0<2>/I0<2>/I0<3>/Q	I0<2>/I0<2>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl234	I0<2>/I0<2>/I0<3>/Q#2	I0<2>/I0<2>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl235	I0<2>/I0<2>/I0<2>/Q	I0<2>/I0<2>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl236	I0<2>/I0<2>/I0<2>/Q#2	I0<2>/I0<2>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl237	I0<2>/I0<2>/I0<1>/Q	I0<2>/I0<2>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl238	I0<2>/I0<2>/I0<1>/Q#2	I0<2>/I0<2>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl239	I0<2>/I0<2>/I0<0>/Q	I0<2>/I0<2>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl240	I0<2>/I0<2>/I0<0>/Q#2	I0<2>/I0<2>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl241	I0<2>/I0<1>/I0<3>/Q	I0<2>/I0<1>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl242	I0<2>/I0<1>/I0<3>/Q#2	I0<2>/I0<1>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl243	I0<2>/I0<1>/I0<2>/Q	I0<2>/I0<1>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl244	I0<2>/I0<1>/I0<2>/Q#2	I0<2>/I0<1>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl245	I0<2>/I0<1>/I0<1>/Q	I0<2>/I0<1>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl246	I0<2>/I0<1>/I0<1>/Q#2	I0<2>/I0<1>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl247	I0<2>/I0<1>/I0<0>/Q	I0<2>/I0<1>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl248	I0<2>/I0<1>/I0<0>/Q#2	I0<2>/I0<1>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl249	I0<2>/I0<0>/I0<3>/Q	I0<2>/I0<0>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl250	I0<2>/I0<0>/I0<3>/Q#2	I0<2>/I0<0>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl251	I0<2>/I0<0>/I0<2>/Q	I0<2>/I0<0>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl252	I0<2>/I0<0>/I0<2>/Q#2	I0<2>/I0<0>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl253	I0<2>/I0<0>/I0<1>/Q	I0<2>/I0<0>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl254	I0<2>/I0<0>/I0<1>/Q#2	I0<2>/I0<0>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl255	I0<2>/I0<0>/I0<0>/Q	I0<2>/I0<0>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl256	I0<2>/I0<0>/I0<0>/Q#2	I0<2>/I0<0>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl257	I0<1>/I0<3>/I0<3>/Q	I0<1>/I0<3>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl258	I0<1>/I0<3>/I0<3>/Q#2	I0<1>/I0<3>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl259	I0<1>/I0<3>/I0<2>/Q	I0<1>/I0<3>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl260	I0<1>/I0<3>/I0<2>/Q#2	I0<1>/I0<3>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl261	I0<1>/I0<3>/I0<1>/Q	I0<1>/I0<3>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl262	I0<1>/I0<3>/I0<1>/Q#2	I0<1>/I0<3>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl263	I0<1>/I0<3>/I0<0>/Q	I0<1>/I0<3>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl264	I0<1>/I0<3>/I0<0>/Q#2	I0<1>/I0<3>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl265	I0<1>/I0<2>/I0<3>/Q	I0<1>/I0<2>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl266	I0<1>/I0<2>/I0<3>/Q#2	I0<1>/I0<2>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl267	I0<1>/I0<2>/I0<2>/Q	I0<1>/I0<2>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl268	I0<1>/I0<2>/I0<2>/Q#2	I0<1>/I0<2>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl269	I0<1>/I0<2>/I0<1>/Q	I0<1>/I0<2>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl270	I0<1>/I0<2>/I0<1>/Q#2	I0<1>/I0<2>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl271	I0<1>/I0<2>/I0<0>/Q	I0<1>/I0<2>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl272	I0<1>/I0<2>/I0<0>/Q#2	I0<1>/I0<2>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl273	I0<1>/I0<1>/I0<3>/Q	I0<1>/I0<1>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl274	I0<1>/I0<1>/I0<3>/Q#2	I0<1>/I0<1>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl275	I0<1>/I0<1>/I0<2>/Q	I0<1>/I0<1>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl276	I0<1>/I0<1>/I0<2>/Q#2	I0<1>/I0<1>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl277	I0<1>/I0<1>/I0<1>/Q	I0<1>/I0<1>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl278	I0<1>/I0<1>/I0<1>/Q#2	I0<1>/I0<1>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl279	I0<1>/I0<1>/I0<0>/Q	I0<1>/I0<1>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl280	I0<1>/I0<1>/I0<0>/Q#2	I0<1>/I0<1>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl281	I0<1>/I0<0>/I0<3>/Q	I0<1>/I0<0>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl282	I0<1>/I0<0>/I0<3>/Q#2	I0<1>/I0<0>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl283	I0<1>/I0<0>/I0<2>/Q	I0<1>/I0<0>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl284	I0<1>/I0<0>/I0<2>/Q#2	I0<1>/I0<0>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl285	I0<1>/I0<0>/I0<1>/Q	I0<1>/I0<0>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl286	I0<1>/I0<0>/I0<1>/Q#2	I0<1>/I0<0>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl287	I0<1>/I0<0>/I0<0>/Q	I0<1>/I0<0>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl288	I0<1>/I0<0>/I0<0>/Q#2	I0<1>/I0<0>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl289	I0<0>/I0<3>/I0<3>/Q	I0<0>/I0<3>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl290	I0<0>/I0<3>/I0<3>/Q#2	I0<0>/I0<3>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl291	I0<0>/I0<3>/I0<2>/Q	I0<0>/I0<3>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl292	I0<0>/I0<3>/I0<2>/Q#2	I0<0>/I0<3>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl293	I0<0>/I0<3>/I0<1>/Q	I0<0>/I0<3>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl294	I0<0>/I0<3>/I0<1>/Q#2	I0<0>/I0<3>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl295	I0<0>/I0<3>/I0<0>/Q	I0<0>/I0<3>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl296	I0<0>/I0<3>/I0<0>/Q#2	I0<0>/I0<3>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl297	I0<0>/I0<2>/I0<3>/Q	I0<0>/I0<2>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl298	I0<0>/I0<2>/I0<3>/Q#2	I0<0>/I0<2>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl299	I0<0>/I0<2>/I0<2>/Q	I0<0>/I0<2>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl300	I0<0>/I0<2>/I0<2>/Q#2	I0<0>/I0<2>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl301	I0<0>/I0<2>/I0<1>/Q	I0<0>/I0<2>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl302	I0<0>/I0<2>/I0<1>/Q#2	I0<0>/I0<2>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl303	I0<0>/I0<2>/I0<0>/Q	I0<0>/I0<2>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl304	I0<0>/I0<2>/I0<0>/Q#2	I0<0>/I0<2>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl305	I0<0>/I0<1>/I0<3>/Q	I0<0>/I0<1>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl306	I0<0>/I0<1>/I0<3>/Q#2	I0<0>/I0<1>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl307	I0<0>/I0<1>/I0<2>/Q	I0<0>/I0<1>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl308	I0<0>/I0<1>/I0<2>/Q#2	I0<0>/I0<1>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl309	I0<0>/I0<1>/I0<1>/Q	I0<0>/I0<1>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl310	I0<0>/I0<1>/I0<1>/Q#2	I0<0>/I0<1>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl311	I0<0>/I0<1>/I0<0>/Q	I0<0>/I0<1>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl312	I0<0>/I0<1>/I0<0>/Q#2	I0<0>/I0<1>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl313	I0<0>/I0<0>/I0<3>/Q	I0<0>/I0<0>/I0<3>/Q#2	   56.4103
+ $poly_conn
Rl314	I0<0>/I0<0>/I0<3>/Q#2	I0<0>/I0<0>/I0<3>/Q#3	   90.3330
+ $poly_conn
Rl315	I0<0>/I0<0>/I0<2>/Q	I0<0>/I0<0>/I0<2>/Q#2	   56.4103
+ $poly_conn
Rl316	I0<0>/I0<0>/I0<2>/Q#2	I0<0>/I0<0>/I0<2>/Q#3	   90.3330
+ $poly_conn
Rl317	I0<0>/I0<0>/I0<1>/Q	I0<0>/I0<0>/I0<1>/Q#2	   56.4103
+ $poly_conn
Rl318	I0<0>/I0<0>/I0<1>/Q#2	I0<0>/I0<0>/I0<1>/Q#3	   90.3330
+ $poly_conn
Rl319	I0<0>/I0<0>/I0<0>/Q	I0<0>/I0<0>/I0<0>/Q#2	   56.4103
+ $poly_conn
Rl320	I0<0>/I0<0>/I0<0>/Q#2	I0<0>/I0<0>/I0<0>/Q#3	   90.3330
+ $poly_conn
Rl321	WL<63>#3	WL<63>#4	  104.7064	$poly_conn
Rl322	WL<62>#3	WL<62>#4	  104.7064	$poly_conn
Rl323	WL<61>#3	WL<61>#4	  104.7064	$poly_conn
Rl324	WL<60>#3	WL<60>#4	  104.7064	$poly_conn
Rl325	WL<59>#3	WL<59>#4	  104.7064	$poly_conn
Rl326	WL<58>#3	WL<58>#4	  104.7064	$poly_conn
Rl327	WL<57>#3	WL<57>#4	  104.7064	$poly_conn
Rl328	WL<56>#3	WL<56>#4	  104.7064	$poly_conn
Rl329	WL<55>#3	WL<55>#4	  104.7064	$poly_conn
Rl330	WL<54>#3	WL<54>#4	  104.7064	$poly_conn
Rl331	WL<53>#3	WL<53>#4	  104.7064	$poly_conn
Rl332	WL<52>#3	WL<52>#4	  104.7064	$poly_conn
Rl333	WL<51>#3	WL<51>#4	  104.7064	$poly_conn
Rl334	WL<50>#3	WL<50>#4	  104.7064	$poly_conn
Rl335	WL<49>#3	WL<49>#4	  104.7064	$poly_conn
Rl336	WL<48>#3	WL<48>#4	  104.7064	$poly_conn
Rl337	WL<47>#3	WL<47>#4	  104.7064	$poly_conn
Rl338	WL<46>#3	WL<46>#4	  104.7064	$poly_conn
Rl339	WL<45>#3	WL<45>#4	  104.7064	$poly_conn
Rl340	WL<44>#3	WL<44>#4	  104.7064	$poly_conn
Rl341	WL<43>#3	WL<43>#4	  104.7064	$poly_conn
Rl342	WL<42>#3	WL<42>#4	  104.7064	$poly_conn
Rl343	WL<41>#3	WL<41>#4	  104.7064	$poly_conn
Rl344	WL<40>#3	WL<40>#4	  104.7064	$poly_conn
Rl345	WL<39>#3	WL<39>#4	  104.7064	$poly_conn
Rl346	WL<38>#3	WL<38>#4	  104.7064	$poly_conn
Rl347	WL<37>#3	WL<37>#4	  104.7064	$poly_conn
Rl348	WL<36>#3	WL<36>#4	  104.7064	$poly_conn
Rl349	WL<35>#3	WL<35>#4	  104.7064	$poly_conn
Rl350	WL<34>#3	WL<34>#4	  104.7064	$poly_conn
Rl351	WL<33>#3	WL<33>#4	  104.7064	$poly_conn
Rl352	WL<32>#3	WL<32>#4	  104.7064	$poly_conn
Rl353	WL<31>#3	WL<31>#4	  104.7064	$poly_conn
Rl354	WL<30>#3	WL<30>#4	  104.7064	$poly_conn
Rl355	WL<29>#3	WL<29>#4	  104.7064	$poly_conn
Rl356	WL<28>#3	WL<28>#4	  104.7064	$poly_conn
Rl357	WL<27>#3	WL<27>#4	  104.7064	$poly_conn
Rl358	WL<26>#3	WL<26>#4	  104.7064	$poly_conn
Rl359	WL<25>#3	WL<25>#4	  104.7064	$poly_conn
Rl360	WL<24>#3	WL<24>#4	  104.7064	$poly_conn
Rl361	WL<23>#3	WL<23>#4	  104.7064	$poly_conn
Rl362	WL<22>#3	WL<22>#4	  104.7064	$poly_conn
Rl363	WL<21>#3	WL<21>#4	  104.7064	$poly_conn
Rl364	WL<20>#3	WL<20>#4	  104.7064	$poly_conn
Rl365	WL<19>#3	WL<19>#4	  104.7064	$poly_conn
Rl366	WL<18>#3	WL<18>#4	  104.7064	$poly_conn
Rl367	WL<17>#3	WL<17>#4	  104.7064	$poly_conn
Rl368	WL<16>#3	WL<16>#4	  104.7064	$poly_conn
Rl369	WL<15>#3	WL<15>#4	  104.7064	$poly_conn
Rl370	WL<14>#3	WL<14>#4	  104.7064	$poly_conn
Rl371	WL<13>#3	WL<13>#4	  104.7064	$poly_conn
Rl372	WL<12>#3	WL<12>#4	  104.7064	$poly_conn
Rl373	WL<11>#3	WL<11>#4	  104.7064	$poly_conn
Rl374	WL<10>#3	WL<10>#4	  104.7064	$poly_conn
Rl375	WL<9>#3	WL<9>#4	  104.7064	$poly_conn
Rl376	WL<8>#3	WL<8>#4	  104.7064	$poly_conn
Rl377	WL<7>#3	WL<7>#4	  104.7064	$poly_conn
Rl378	WL<6>#3	WL<6>#4	  104.7064	$poly_conn
Rl379	WL<5>#3	WL<5>#4	  104.7064	$poly_conn
Rl380	WL<4>#3	WL<4>#4	  104.7064	$poly_conn
Rl381	WL<3>#3	WL<3>#4	  104.7064	$poly_conn
Rl382	WL<2>#3	WL<2>#4	  104.7064	$poly_conn
Rl383	WL<1>#3	WL<1>#4	  104.7064	$poly_conn
Rl384	WL<0>#3	WL<0>#4	  104.7064	$poly_conn
Rk1	WL<63>#2	WL<63>#5	    6.6000	$metal1_conn
Rk2	WL<62>#2	WL<62>#5	    6.6000	$metal1_conn
Rk3	WL<61>#2	WL<61>#5	    6.6000	$metal1_conn
Rk4	WL<60>#2	WL<60>#5	    6.6000	$metal1_conn
Rk5	WL<59>#2	WL<59>#5	    6.6000	$metal1_conn
Rk6	WL<58>#2	WL<58>#5	    6.6000	$metal1_conn
Rk7	WL<57>#2	WL<57>#5	    6.6000	$metal1_conn
Rk8	WL<56>#2	WL<56>#5	    6.6000	$metal1_conn
Rk9	WL<55>#2	WL<55>#5	    6.6000	$metal1_conn
Rk10	WL<54>#2	WL<54>#5	    6.6000	$metal1_conn
Rk11	WL<53>#2	WL<53>#5	    6.6000	$metal1_conn
Rk12	WL<52>#2	WL<52>#5	    6.6000	$metal1_conn
Rk13	WL<51>#2	WL<51>#5	    6.6000	$metal1_conn
Rk14	WL<50>#2	WL<50>#5	    6.6000	$metal1_conn
Rk15	WL<49>#2	WL<49>#5	    6.6000	$metal1_conn
Rk16	WL<48>#2	WL<48>#5	    6.6000	$metal1_conn
Rk17	WL<47>#2	WL<47>#5	    6.6000	$metal1_conn
Rk18	WL<46>#2	WL<46>#5	    6.6000	$metal1_conn
Rk19	WL<45>#2	WL<45>#5	    6.6000	$metal1_conn
Rk20	WL<44>#2	WL<44>#5	    6.6000	$metal1_conn
Rk21	WL<43>#2	WL<43>#5	    6.6000	$metal1_conn
Rk22	WL<42>#2	WL<42>#5	    6.6000	$metal1_conn
Rk23	WL<41>#2	WL<41>#5	    6.6000	$metal1_conn
Rk24	WL<40>#2	WL<40>#5	    6.6000	$metal1_conn
Rk25	WL<39>#2	WL<39>#5	    6.6000	$metal1_conn
Rk26	WL<38>#2	WL<38>#5	    6.6000	$metal1_conn
Rk27	WL<37>#2	WL<37>#5	    6.6000	$metal1_conn
Rk28	WL<36>#2	WL<36>#5	    6.6000	$metal1_conn
Rk29	WL<35>#2	WL<35>#5	    6.6000	$metal1_conn
Rk30	WL<34>#2	WL<34>#5	    6.6000	$metal1_conn
Rk31	WL<33>#2	WL<33>#5	    6.6000	$metal1_conn
Rk32	WL<32>#2	WL<32>#5	    6.6000	$metal1_conn
Rk33	WL<31>#2	WL<31>#5	    6.6000	$metal1_conn
Rk34	WL<30>#2	WL<30>#5	    6.6000	$metal1_conn
Rk35	WL<29>#2	WL<29>#5	    6.6000	$metal1_conn
Rk36	WL<28>#2	WL<28>#5	    6.6000	$metal1_conn
Rk37	WL<27>#2	WL<27>#5	    6.6000	$metal1_conn
Rk38	WL<26>#2	WL<26>#5	    6.6000	$metal1_conn
Rk39	WL<25>#2	WL<25>#5	    6.6000	$metal1_conn
Rk40	WL<24>#2	WL<24>#5	    6.6000	$metal1_conn
Rk41	WL<23>#2	WL<23>#5	    6.6000	$metal1_conn
Rk42	WL<22>#2	WL<22>#5	    6.6000	$metal1_conn
Rk43	WL<21>#2	WL<21>#5	    6.6000	$metal1_conn
Rk44	WL<20>#2	WL<20>#5	    6.6000	$metal1_conn
Rk45	WL<19>#2	WL<19>#5	    6.6000	$metal1_conn
Rk46	WL<18>#2	WL<18>#5	    6.6000	$metal1_conn
Rk47	WL<17>#2	WL<17>#5	    6.6000	$metal1_conn
Rk48	WL<16>#2	WL<16>#5	    6.6000	$metal1_conn
Rk49	WL<15>#2	WL<15>#5	    6.6000	$metal1_conn
Rk50	WL<14>#2	WL<14>#5	    6.6000	$metal1_conn
Rk51	WL<13>#2	WL<13>#5	    6.6000	$metal1_conn
Rk52	WL<12>#2	WL<12>#5	    6.6000	$metal1_conn
Rk53	WL<11>#2	WL<11>#5	    6.6000	$metal1_conn
Rk54	WL<10>#2	WL<10>#5	    6.6000	$metal1_conn
Rk55	WL<9>#2	WL<9>#5	    6.6000	$metal1_conn
Rk56	WL<8>#2	WL<8>#5	    6.6000	$metal1_conn
Rk57	WL<7>#2	WL<7>#5	    6.6000	$metal1_conn
Rk58	WL<6>#2	WL<6>#5	    6.6000	$metal1_conn
Rk59	WL<5>#2	WL<5>#5	    6.6000	$metal1_conn
Rk60	WL<4>#2	WL<4>#5	    6.6000	$metal1_conn
Rk61	WL<3>#2	WL<3>#5	    6.6000	$metal1_conn
Rk62	WL<2>#2	WL<2>#5	    6.6000	$metal1_conn
Rk63	WL<1>#2	WL<1>#5	    6.6000	$metal1_conn
Rk64	WL<0>#2	WL<0>#5	    6.6000	$metal1_conn
Rk65	VSS#1	VSS#2	   27.3722	$metal1_conn
Rk66	VSS#1	VSS#3	   27.3722	$metal1_conn
Rk67	VSS#4	VSS#5	   81.7666	$metal1_conn
Rk68	VSS#6	VSS#7	   81.7666	$metal1_conn
Rk69	VSS#8	VSS#9	   81.7666	$metal1_conn
Rk70	VSS#10	VSS#11	   81.7666	$metal1_conn
Rk71	VSS#12	VSS#13	   81.7666	$metal1_conn
Rk72	VSS#14	VSS#15	   81.7666	$metal1_conn
Rk73	VSS#16	VSS#17	   81.7666	$metal1_conn
Rk74	VSS#18	VSS#19	   81.7666	$metal1_conn
Rk75	VSS#20	VSS#21	   81.7666	$metal1_conn
Rk76	VSS#22	VSS#23	   81.7666	$metal1_conn
Rk77	VSS#24	VSS#25	   81.7666	$metal1_conn
Rk78	VSS#26	VSS#27	   81.7666	$metal1_conn
Rk79	VSS#28	VSS#29	   81.7666	$metal1_conn
Rk80	VSS#30	VSS#31	   81.7666	$metal1_conn
Rk81	VSS#32	VSS#33	   81.7666	$metal1_conn
Rk82	VSS#34	VSS#35	   81.7666	$metal1_conn
Rk83	VSS#36	VSS#37	   81.7666	$metal1_conn
Rk84	VSS#38	VSS#39	   81.7666	$metal1_conn
Rk85	VSS#40	VSS#41	   81.7666	$metal1_conn
Rk86	VSS#42	VSS#43	   81.7666	$metal1_conn
Rk87	VSS#44	VSS#45	   81.7666	$metal1_conn
Rk88	VSS#46	VSS#47	   81.7666	$metal1_conn
Rk89	VSS#48	VSS#49	   81.7666	$metal1_conn
Rk90	VSS#50	VSS#51	   81.7666	$metal1_conn
Rk91	VSS#52	VSS#53	   81.7666	$metal1_conn
Rk92	VSS#54	VSS#55	   81.7666	$metal1_conn
Rk93	VSS#56	VSS#57	   81.7666	$metal1_conn
Rk94	VSS#58	VSS#59	   81.7666	$metal1_conn
Rk95	VSS#60	VSS#61	   81.7666	$metal1_conn
Rk96	VSS#62	VSS#63	   81.7666	$metal1_conn
Rk97	VSS#64	VSS#65	   81.7666	$metal1_conn
Rk98	VSS#66	VSS#67	   81.7666	$metal1_conn
Rk99	VSS#68	VSS#69	   81.7666	$metal1_conn
Rk100	BL#1	BL#2	   81.6000	$metal1_conn
Rk101	BL#3	BL#4	   81.6000	$metal1_conn
Rk102	BL#5	BL#6	   81.6000	$metal1_conn
Rk103	BL#7	BL#8	   81.6000	$metal1_conn
Rk104	BL#9	BL#10	   81.6000	$metal1_conn
Rk105	BL#11	BL#12	   81.6000	$metal1_conn
Rk106	BL#13	BL#14	   81.6000	$metal1_conn
Rk107	BL#15	BL#16	   81.6000	$metal1_conn
Rk108	BL#17	BL#18	   81.6000	$metal1_conn
Rk109	BL#19	BL#20	   81.6000	$metal1_conn
Rk110	BL#21	BL#22	   81.6000	$metal1_conn
Rk111	BL#23	BL#24	   81.6000	$metal1_conn
Rk112	BL#25	BL#26	   81.6000	$metal1_conn
Rk113	BL#27	BL#28	   81.6000	$metal1_conn
Rk114	BL#29	BL#30	   81.6000	$metal1_conn
Rk115	BL#31	BL#32	   81.6000	$metal1_conn
Rk116	BL#33	BL#34	   81.6000	$metal1_conn
Rk117	BL#35	BL#36	   81.6000	$metal1_conn
Rk118	BL#37	BL#38	   81.6000	$metal1_conn
Rk119	BL#39	BL#40	   81.6000	$metal1_conn
Rk120	BL#41	BL#42	   81.6000	$metal1_conn
Rk121	BL#43	BL#44	   81.6000	$metal1_conn
Rk122	BL#45	BL#46	   81.6000	$metal1_conn
Rk123	BL#47	BL#48	   81.6000	$metal1_conn
Rk124	BL#49	BL#50	   81.6000	$metal1_conn
Rk125	BL#51	BL#52	   81.6000	$metal1_conn
Rk126	BL#53	BL#54	   81.6000	$metal1_conn
Rk127	BL#55	BL#56	   81.6000	$metal1_conn
Rk128	BL#57	BL#58	   81.6000	$metal1_conn
Rk129	BL#59	BL#60	   81.6000	$metal1_conn
Rk130	BL#61	BL#62	   81.6000	$metal1_conn
Rk131	BL#63	BL#64	   81.6000	$metal1_conn
Rk132	I0<3>/I0<3>/I0<3>/Q#3	I0<3>/I0<3>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk133	I0<3>/I0<3>/I0<3>/Q#5	I0<3>/I0<3>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk134	I0<3>/I0<3>/I0<3>/Q#4	I0<3>/I0<3>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk135	I0<3>/I0<3>/I0<2>/Q#3	I0<3>/I0<3>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk136	I0<3>/I0<3>/I0<2>/Q#5	I0<3>/I0<3>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk137	I0<3>/I0<3>/I0<2>/Q#4	I0<3>/I0<3>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk138	I0<3>/I0<3>/I0<1>/Q#3	I0<3>/I0<3>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk139	I0<3>/I0<3>/I0<1>/Q#5	I0<3>/I0<3>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk140	I0<3>/I0<3>/I0<1>/Q#4	I0<3>/I0<3>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk141	I0<3>/I0<3>/I0<0>/Q#3	I0<3>/I0<3>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk142	I0<3>/I0<3>/I0<0>/Q#5	I0<3>/I0<3>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk143	I0<3>/I0<3>/I0<0>/Q#4	I0<3>/I0<3>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk144	I0<3>/I0<2>/I0<3>/Q#3	I0<3>/I0<2>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk145	I0<3>/I0<2>/I0<3>/Q#5	I0<3>/I0<2>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk146	I0<3>/I0<2>/I0<3>/Q#4	I0<3>/I0<2>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk147	I0<3>/I0<2>/I0<2>/Q#3	I0<3>/I0<2>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk148	I0<3>/I0<2>/I0<2>/Q#5	I0<3>/I0<2>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk149	I0<3>/I0<2>/I0<2>/Q#4	I0<3>/I0<2>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk150	I0<3>/I0<2>/I0<1>/Q#3	I0<3>/I0<2>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk151	I0<3>/I0<2>/I0<1>/Q#5	I0<3>/I0<2>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk152	I0<3>/I0<2>/I0<1>/Q#4	I0<3>/I0<2>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk153	I0<3>/I0<2>/I0<0>/Q#3	I0<3>/I0<2>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk154	I0<3>/I0<2>/I0<0>/Q#5	I0<3>/I0<2>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk155	I0<3>/I0<2>/I0<0>/Q#4	I0<3>/I0<2>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk156	I0<3>/I0<1>/I0<3>/Q#3	I0<3>/I0<1>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk157	I0<3>/I0<1>/I0<3>/Q#5	I0<3>/I0<1>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk158	I0<3>/I0<1>/I0<3>/Q#4	I0<3>/I0<1>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk159	I0<3>/I0<1>/I0<2>/Q#3	I0<3>/I0<1>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk160	I0<3>/I0<1>/I0<2>/Q#5	I0<3>/I0<1>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk161	I0<3>/I0<1>/I0<2>/Q#4	I0<3>/I0<1>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk162	I0<3>/I0<1>/I0<1>/Q#3	I0<3>/I0<1>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk163	I0<3>/I0<1>/I0<1>/Q#5	I0<3>/I0<1>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk164	I0<3>/I0<1>/I0<1>/Q#4	I0<3>/I0<1>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk165	I0<3>/I0<1>/I0<0>/Q#3	I0<3>/I0<1>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk166	I0<3>/I0<1>/I0<0>/Q#5	I0<3>/I0<1>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk167	I0<3>/I0<1>/I0<0>/Q#4	I0<3>/I0<1>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk168	I0<3>/I0<0>/I0<3>/Q#3	I0<3>/I0<0>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk169	I0<3>/I0<0>/I0<3>/Q#5	I0<3>/I0<0>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk170	I0<3>/I0<0>/I0<3>/Q#4	I0<3>/I0<0>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk171	I0<3>/I0<0>/I0<2>/Q#3	I0<3>/I0<0>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk172	I0<3>/I0<0>/I0<2>/Q#5	I0<3>/I0<0>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk173	I0<3>/I0<0>/I0<2>/Q#4	I0<3>/I0<0>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk174	I0<3>/I0<0>/I0<1>/Q#3	I0<3>/I0<0>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk175	I0<3>/I0<0>/I0<1>/Q#5	I0<3>/I0<0>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk176	I0<3>/I0<0>/I0<1>/Q#4	I0<3>/I0<0>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk177	I0<3>/I0<0>/I0<0>/Q#3	I0<3>/I0<0>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk178	I0<3>/I0<0>/I0<0>/Q#5	I0<3>/I0<0>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk179	I0<3>/I0<0>/I0<0>/Q#4	I0<3>/I0<0>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk180	I0<2>/I0<3>/I0<3>/Q#3	I0<2>/I0<3>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk181	I0<2>/I0<3>/I0<3>/Q#5	I0<2>/I0<3>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk182	I0<2>/I0<3>/I0<3>/Q#4	I0<2>/I0<3>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk183	I0<2>/I0<3>/I0<2>/Q#3	I0<2>/I0<3>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk184	I0<2>/I0<3>/I0<2>/Q#5	I0<2>/I0<3>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk185	I0<2>/I0<3>/I0<2>/Q#4	I0<2>/I0<3>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk186	I0<2>/I0<3>/I0<1>/Q#3	I0<2>/I0<3>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk187	I0<2>/I0<3>/I0<1>/Q#5	I0<2>/I0<3>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk188	I0<2>/I0<3>/I0<1>/Q#4	I0<2>/I0<3>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk189	I0<2>/I0<3>/I0<0>/Q#3	I0<2>/I0<3>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk190	I0<2>/I0<3>/I0<0>/Q#5	I0<2>/I0<3>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk191	I0<2>/I0<3>/I0<0>/Q#4	I0<2>/I0<3>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk192	I0<2>/I0<2>/I0<3>/Q#3	I0<2>/I0<2>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk193	I0<2>/I0<2>/I0<3>/Q#5	I0<2>/I0<2>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk194	I0<2>/I0<2>/I0<3>/Q#4	I0<2>/I0<2>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk195	I0<2>/I0<2>/I0<2>/Q#3	I0<2>/I0<2>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk196	I0<2>/I0<2>/I0<2>/Q#5	I0<2>/I0<2>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk197	I0<2>/I0<2>/I0<2>/Q#4	I0<2>/I0<2>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk198	I0<2>/I0<2>/I0<1>/Q#3	I0<2>/I0<2>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk199	I0<2>/I0<2>/I0<1>/Q#5	I0<2>/I0<2>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk200	I0<2>/I0<2>/I0<1>/Q#4	I0<2>/I0<2>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk201	I0<2>/I0<2>/I0<0>/Q#3	I0<2>/I0<2>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk202	I0<2>/I0<2>/I0<0>/Q#5	I0<2>/I0<2>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk203	I0<2>/I0<2>/I0<0>/Q#4	I0<2>/I0<2>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk204	I0<2>/I0<1>/I0<3>/Q#3	I0<2>/I0<1>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk205	I0<2>/I0<1>/I0<3>/Q#5	I0<2>/I0<1>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk206	I0<2>/I0<1>/I0<3>/Q#4	I0<2>/I0<1>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk207	I0<2>/I0<1>/I0<2>/Q#3	I0<2>/I0<1>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk208	I0<2>/I0<1>/I0<2>/Q#5	I0<2>/I0<1>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk209	I0<2>/I0<1>/I0<2>/Q#4	I0<2>/I0<1>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk210	I0<2>/I0<1>/I0<1>/Q#3	I0<2>/I0<1>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk211	I0<2>/I0<1>/I0<1>/Q#5	I0<2>/I0<1>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk212	I0<2>/I0<1>/I0<1>/Q#4	I0<2>/I0<1>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk213	I0<2>/I0<1>/I0<0>/Q#3	I0<2>/I0<1>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk214	I0<2>/I0<1>/I0<0>/Q#5	I0<2>/I0<1>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk215	I0<2>/I0<1>/I0<0>/Q#4	I0<2>/I0<1>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk216	I0<2>/I0<0>/I0<3>/Q#3	I0<2>/I0<0>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk217	I0<2>/I0<0>/I0<3>/Q#5	I0<2>/I0<0>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk218	I0<2>/I0<0>/I0<3>/Q#4	I0<2>/I0<0>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk219	I0<2>/I0<0>/I0<2>/Q#3	I0<2>/I0<0>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk220	I0<2>/I0<0>/I0<2>/Q#5	I0<2>/I0<0>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk221	I0<2>/I0<0>/I0<2>/Q#4	I0<2>/I0<0>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk222	I0<2>/I0<0>/I0<1>/Q#3	I0<2>/I0<0>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk223	I0<2>/I0<0>/I0<1>/Q#5	I0<2>/I0<0>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk224	I0<2>/I0<0>/I0<1>/Q#4	I0<2>/I0<0>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk225	I0<2>/I0<0>/I0<0>/Q#3	I0<2>/I0<0>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk226	I0<2>/I0<0>/I0<0>/Q#5	I0<2>/I0<0>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk227	I0<2>/I0<0>/I0<0>/Q#4	I0<2>/I0<0>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk228	I0<1>/I0<3>/I0<3>/Q#3	I0<1>/I0<3>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk229	I0<1>/I0<3>/I0<3>/Q#5	I0<1>/I0<3>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk230	I0<1>/I0<3>/I0<3>/Q#4	I0<1>/I0<3>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk231	I0<1>/I0<3>/I0<2>/Q#3	I0<1>/I0<3>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk232	I0<1>/I0<3>/I0<2>/Q#5	I0<1>/I0<3>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk233	I0<1>/I0<3>/I0<2>/Q#4	I0<1>/I0<3>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk234	I0<1>/I0<3>/I0<1>/Q#3	I0<1>/I0<3>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk235	I0<1>/I0<3>/I0<1>/Q#5	I0<1>/I0<3>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk236	I0<1>/I0<3>/I0<1>/Q#4	I0<1>/I0<3>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk237	I0<1>/I0<3>/I0<0>/Q#3	I0<1>/I0<3>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk238	I0<1>/I0<3>/I0<0>/Q#5	I0<1>/I0<3>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk239	I0<1>/I0<3>/I0<0>/Q#4	I0<1>/I0<3>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk240	I0<1>/I0<2>/I0<3>/Q#3	I0<1>/I0<2>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk241	I0<1>/I0<2>/I0<3>/Q#5	I0<1>/I0<2>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk242	I0<1>/I0<2>/I0<3>/Q#4	I0<1>/I0<2>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk243	I0<1>/I0<2>/I0<2>/Q#3	I0<1>/I0<2>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk244	I0<1>/I0<2>/I0<2>/Q#5	I0<1>/I0<2>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk245	I0<1>/I0<2>/I0<2>/Q#4	I0<1>/I0<2>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk246	I0<1>/I0<2>/I0<1>/Q#3	I0<1>/I0<2>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk247	I0<1>/I0<2>/I0<1>/Q#5	I0<1>/I0<2>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk248	I0<1>/I0<2>/I0<1>/Q#4	I0<1>/I0<2>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk249	I0<1>/I0<2>/I0<0>/Q#3	I0<1>/I0<2>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk250	I0<1>/I0<2>/I0<0>/Q#5	I0<1>/I0<2>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk251	I0<1>/I0<2>/I0<0>/Q#4	I0<1>/I0<2>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk252	I0<1>/I0<1>/I0<3>/Q#3	I0<1>/I0<1>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk253	I0<1>/I0<1>/I0<3>/Q#5	I0<1>/I0<1>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk254	I0<1>/I0<1>/I0<3>/Q#4	I0<1>/I0<1>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk255	I0<1>/I0<1>/I0<2>/Q#3	I0<1>/I0<1>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk256	I0<1>/I0<1>/I0<2>/Q#5	I0<1>/I0<1>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk257	I0<1>/I0<1>/I0<2>/Q#4	I0<1>/I0<1>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk258	I0<1>/I0<1>/I0<1>/Q#3	I0<1>/I0<1>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk259	I0<1>/I0<1>/I0<1>/Q#5	I0<1>/I0<1>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk260	I0<1>/I0<1>/I0<1>/Q#4	I0<1>/I0<1>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk261	I0<1>/I0<1>/I0<0>/Q#3	I0<1>/I0<1>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk262	I0<1>/I0<1>/I0<0>/Q#5	I0<1>/I0<1>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk263	I0<1>/I0<1>/I0<0>/Q#4	I0<1>/I0<1>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk264	I0<1>/I0<0>/I0<3>/Q#3	I0<1>/I0<0>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk265	I0<1>/I0<0>/I0<3>/Q#5	I0<1>/I0<0>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk266	I0<1>/I0<0>/I0<3>/Q#4	I0<1>/I0<0>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk267	I0<1>/I0<0>/I0<2>/Q#3	I0<1>/I0<0>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk268	I0<1>/I0<0>/I0<2>/Q#5	I0<1>/I0<0>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk269	I0<1>/I0<0>/I0<2>/Q#4	I0<1>/I0<0>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk270	I0<1>/I0<0>/I0<1>/Q#3	I0<1>/I0<0>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk271	I0<1>/I0<0>/I0<1>/Q#5	I0<1>/I0<0>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk272	I0<1>/I0<0>/I0<1>/Q#4	I0<1>/I0<0>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk273	I0<1>/I0<0>/I0<0>/Q#3	I0<1>/I0<0>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk274	I0<1>/I0<0>/I0<0>/Q#5	I0<1>/I0<0>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk275	I0<1>/I0<0>/I0<0>/Q#4	I0<1>/I0<0>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk276	I0<0>/I0<3>/I0<3>/Q#3	I0<0>/I0<3>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk277	I0<0>/I0<3>/I0<3>/Q#5	I0<0>/I0<3>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk278	I0<0>/I0<3>/I0<3>/Q#4	I0<0>/I0<3>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk279	I0<0>/I0<3>/I0<2>/Q#3	I0<0>/I0<3>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk280	I0<0>/I0<3>/I0<2>/Q#5	I0<0>/I0<3>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk281	I0<0>/I0<3>/I0<2>/Q#4	I0<0>/I0<3>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk282	I0<0>/I0<3>/I0<1>/Q#3	I0<0>/I0<3>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk283	I0<0>/I0<3>/I0<1>/Q#5	I0<0>/I0<3>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk284	I0<0>/I0<3>/I0<1>/Q#4	I0<0>/I0<3>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk285	I0<0>/I0<3>/I0<0>/Q#3	I0<0>/I0<3>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk286	I0<0>/I0<3>/I0<0>/Q#5	I0<0>/I0<3>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk287	I0<0>/I0<3>/I0<0>/Q#4	I0<0>/I0<3>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk288	I0<0>/I0<2>/I0<3>/Q#3	I0<0>/I0<2>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk289	I0<0>/I0<2>/I0<3>/Q#5	I0<0>/I0<2>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk290	I0<0>/I0<2>/I0<3>/Q#4	I0<0>/I0<2>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk291	I0<0>/I0<2>/I0<2>/Q#3	I0<0>/I0<2>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk292	I0<0>/I0<2>/I0<2>/Q#5	I0<0>/I0<2>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk293	I0<0>/I0<2>/I0<2>/Q#4	I0<0>/I0<2>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk294	I0<0>/I0<2>/I0<1>/Q#3	I0<0>/I0<2>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk295	I0<0>/I0<2>/I0<1>/Q#5	I0<0>/I0<2>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk296	I0<0>/I0<2>/I0<1>/Q#4	I0<0>/I0<2>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk297	I0<0>/I0<2>/I0<0>/Q#3	I0<0>/I0<2>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk298	I0<0>/I0<2>/I0<0>/Q#5	I0<0>/I0<2>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk299	I0<0>/I0<2>/I0<0>/Q#4	I0<0>/I0<2>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk300	I0<0>/I0<1>/I0<3>/Q#3	I0<0>/I0<1>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk301	I0<0>/I0<1>/I0<3>/Q#5	I0<0>/I0<1>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk302	I0<0>/I0<1>/I0<3>/Q#4	I0<0>/I0<1>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk303	I0<0>/I0<1>/I0<2>/Q#3	I0<0>/I0<1>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk304	I0<0>/I0<1>/I0<2>/Q#5	I0<0>/I0<1>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk305	I0<0>/I0<1>/I0<2>/Q#4	I0<0>/I0<1>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk306	I0<0>/I0<1>/I0<1>/Q#3	I0<0>/I0<1>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk307	I0<0>/I0<1>/I0<1>/Q#5	I0<0>/I0<1>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk308	I0<0>/I0<1>/I0<1>/Q#4	I0<0>/I0<1>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk309	I0<0>/I0<1>/I0<0>/Q#3	I0<0>/I0<1>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk310	I0<0>/I0<1>/I0<0>/Q#5	I0<0>/I0<1>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk311	I0<0>/I0<1>/I0<0>/Q#4	I0<0>/I0<1>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk312	I0<0>/I0<0>/I0<3>/Q#3	I0<0>/I0<0>/I0<3>/Q#5	    0.1682
+ $metal1_conn
Rk313	I0<0>/I0<0>/I0<3>/Q#5	I0<0>/I0<0>/I0<3>/Q#6	   75.2888
+ $metal1_conn
Rk314	I0<0>/I0<0>/I0<3>/Q#4	I0<0>/I0<0>/I0<3>/Q#5	   62.0000
+ $metal1_conn
Rk315	I0<0>/I0<0>/I0<2>/Q#3	I0<0>/I0<0>/I0<2>/Q#5	    0.1682
+ $metal1_conn
Rk316	I0<0>/I0<0>/I0<2>/Q#5	I0<0>/I0<0>/I0<2>/Q#6	   75.2888
+ $metal1_conn
Rk317	I0<0>/I0<0>/I0<2>/Q#4	I0<0>/I0<0>/I0<2>/Q#5	   62.0000
+ $metal1_conn
Rk318	I0<0>/I0<0>/I0<1>/Q#3	I0<0>/I0<0>/I0<1>/Q#5	    0.1682
+ $metal1_conn
Rk319	I0<0>/I0<0>/I0<1>/Q#5	I0<0>/I0<0>/I0<1>/Q#6	   75.2888
+ $metal1_conn
Rk320	I0<0>/I0<0>/I0<1>/Q#4	I0<0>/I0<0>/I0<1>/Q#5	   62.0000
+ $metal1_conn
Rk321	I0<0>/I0<0>/I0<0>/Q#3	I0<0>/I0<0>/I0<0>/Q#5	    0.1682
+ $metal1_conn
Rk322	I0<0>/I0<0>/I0<0>/Q#5	I0<0>/I0<0>/I0<0>/Q#6	   75.2888
+ $metal1_conn
Rk323	I0<0>/I0<0>/I0<0>/Q#4	I0<0>/I0<0>/I0<0>/Q#5	   62.0000
+ $metal1_conn
Rk324	VDD#1	VDD#2	   68.7316	$metal1_conn
Rk325	VDD#3	VDD#4	   68.7324	$metal1_conn
Rk326	VDD#5	VDD#6	   68.7324	$metal1_conn
Rk327	VDD#7	VDD#8	   68.7324	$metal1_conn
Rk328	VDD#9	VDD#10	   68.7324	$metal1_conn
Rk329	VDD#11	VDD#12	   68.7324	$metal1_conn
Rk330	VDD#13	VDD#14	   68.7324	$metal1_conn
Rk331	VDD#15	VDD#16	   68.7324	$metal1_conn
Rk332	VDD#17	VDD#18	   68.7324	$metal1_conn
Rk333	VDD#19	VDD#20	   68.7324	$metal1_conn
Rk334	VDD#21	VDD#22	   68.7324	$metal1_conn
Rk335	VDD#23	VDD#24	   68.7324	$metal1_conn
Rk336	VDD#25	VDD#26	   68.7324	$metal1_conn
Rk337	VDD#27	VDD#28	   68.7324	$metal1_conn
Rk338	VDD#29	VDD#30	   68.7324	$metal1_conn
Rk339	VDD#31	VDD#32	   68.7324	$metal1_conn
Rk340	VDD#33	VDD#34	   68.7324	$metal1_conn
Rk341	VDD#35	VDD#36	   68.7324	$metal1_conn
Rk342	VDD#37	VDD#38	   68.7324	$metal1_conn
Rk343	VDD#39	VDD#40	   68.7324	$metal1_conn
Rk344	VDD#41	VDD#42	   68.7324	$metal1_conn
Rk345	VDD#43	VDD#44	   68.7324	$metal1_conn
Rk346	VDD#45	VDD#46	   68.7324	$metal1_conn
Rk347	VDD#47	VDD#48	   68.7324	$metal1_conn
Rk348	VDD#49	VDD#50	   68.7324	$metal1_conn
Rk349	VDD#51	VDD#52	   68.7324	$metal1_conn
Rk350	VDD#53	VDD#54	   68.7324	$metal1_conn
Rk351	VDD#55	VDD#56	   68.7324	$metal1_conn
Rk352	VDD#57	VDD#58	   68.7324	$metal1_conn
Rk353	VDD#59	VDD#60	   68.7324	$metal1_conn
Rk354	VDD#61	VDD#62	   68.7324	$metal1_conn
Rk355	VDD#63	VDD#64	   68.7324	$metal1_conn
Rk356	VDD#65	VDD#66	   68.7316	$metal1_conn
Rk357	VDD#67	VDD#68	   31.6000	$metal1_conn
Rk358	VDD#69	VDD#68	   31.6000	$metal1_conn
Rk359	VDD#70	VDD#71	   68.7324	$metal1_conn
Rk360	VDD#72	VDD#73	   68.7324	$metal1_conn
Rk361	VDD#74	VDD#75	   68.7324	$metal1_conn
Rk362	VDD#76	VDD#77	   68.7324	$metal1_conn
Rk363	VDD#78	VDD#79	   68.7324	$metal1_conn
Rk364	VDD#80	VDD#81	   68.7324	$metal1_conn
Rk365	VDD#82	VDD#83	   68.7324	$metal1_conn
Rk366	VDD#84	VDD#85	   68.7324	$metal1_conn
Rk367	VDD#86	VDD#87	   68.7324	$metal1_conn
Rk368	VDD#88	VDD#89	   68.7324	$metal1_conn
Rk369	VDD#90	VDD#91	   68.7324	$metal1_conn
Rk370	VDD#92	VDD#93	   68.7324	$metal1_conn
Rk371	VDD#94	VDD#95	   68.7324	$metal1_conn
Rk372	VDD#96	VDD#97	   68.7324	$metal1_conn
Rk373	VDD#98	VDD#99	   68.7324	$metal1_conn
Rk374	VDD#100	VDD#101	   68.7324	$metal1_conn
Rk375	VDD#102	VDD#103	   68.7324	$metal1_conn
Rk376	VDD#104	VDD#105	   68.7324	$metal1_conn
Rk377	VDD#106	VDD#107	   68.7324	$metal1_conn
Rk378	VDD#108	VDD#109	   68.7324	$metal1_conn
Rk379	VDD#110	VDD#111	   68.7324	$metal1_conn
Rk380	VDD#112	VDD#113	   68.7324	$metal1_conn
Rk381	VDD#114	VDD#115	   68.7324	$metal1_conn
Rk382	VDD#116	VDD#117	   68.7324	$metal1_conn
Rk383	VDD#118	VDD#119	   68.7324	$metal1_conn
Rk384	VDD#120	VDD#121	   68.7324	$metal1_conn
Rk385	VDD#122	VDD#123	   68.7324	$metal1_conn
Rk386	VDD#124	VDD#125	   68.7324	$metal1_conn
Rk387	VDD#126	VDD#127	   68.7324	$metal1_conn
Rk388	VDD#128	VDD#129	   68.7324	$metal1_conn
Rk389	VDD#130	VDD#131	   68.7324	$metal1_conn
Rk390	VDD#132	VDD#133	   68.7324	$metal1_conn
Rk391	BLB#1	BLB#2	   81.6000	$metal1_conn
Rk392	BLB#3	BLB#4	   81.6000	$metal1_conn
Rk393	BLB#5	BLB#6	   81.6000	$metal1_conn
Rk394	BLB#7	BLB#8	   81.6000	$metal1_conn
Rk395	BLB#9	BLB#10	   81.6000	$metal1_conn
Rk396	BLB#11	BLB#12	   81.6000	$metal1_conn
Rk397	BLB#13	BLB#14	   81.6000	$metal1_conn
Rk398	BLB#15	BLB#16	   81.6000	$metal1_conn
Rk399	BLB#17	BLB#18	   81.6000	$metal1_conn
Rk400	BLB#19	BLB#20	   81.6000	$metal1_conn
Rk401	BLB#21	BLB#22	   81.6000	$metal1_conn
Rk402	BLB#23	BLB#24	   81.6000	$metal1_conn
Rk403	BLB#25	BLB#26	   81.6000	$metal1_conn
Rk404	BLB#27	BLB#28	   81.6000	$metal1_conn
Rk405	BLB#29	BLB#30	   81.6000	$metal1_conn
Rk406	BLB#31	BLB#32	   81.6000	$metal1_conn
Rk407	BLB#33	BLB#34	   81.6000	$metal1_conn
Rk408	BLB#35	BLB#36	   81.6000	$metal1_conn
Rk409	BLB#37	BLB#38	   81.6000	$metal1_conn
Rk410	BLB#39	BLB#40	   81.6000	$metal1_conn
Rk411	BLB#41	BLB#42	   81.6000	$metal1_conn
Rk412	BLB#43	BLB#44	   81.6000	$metal1_conn
Rk413	BLB#45	BLB#46	   81.6000	$metal1_conn
Rk414	BLB#47	BLB#48	   81.6000	$metal1_conn
Rk415	BLB#49	BLB#50	   81.6000	$metal1_conn
Rk416	BLB#51	BLB#52	   81.6000	$metal1_conn
Rk417	BLB#53	BLB#54	   81.6000	$metal1_conn
Rk418	BLB#55	BLB#56	   81.6000	$metal1_conn
Rk419	BLB#57	BLB#58	   81.6000	$metal1_conn
Rk420	BLB#59	BLB#60	   81.6000	$metal1_conn
Rk421	BLB#61	BLB#62	   81.6000	$metal1_conn
Rk422	BLB#63	BLB#64	   81.6000	$metal1_conn
Rk423	BLB#65	BLB#66	   81.6000	$metal1_conn
Rk424	I0<3>/I0<3>/I0<3>/QB#4	I0<3>/I0<3>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk425	I0<3>/I0<3>/I0<3>/QB#6	I0<3>/I0<3>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk426	I0<3>/I0<3>/I0<3>/QB#5	I0<3>/I0<3>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk427	I0<3>/I0<3>/I0<2>/QB#4	I0<3>/I0<3>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk428	I0<3>/I0<3>/I0<2>/QB#6	I0<3>/I0<3>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk429	I0<3>/I0<3>/I0<2>/QB#5	I0<3>/I0<3>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk430	I0<3>/I0<3>/I0<1>/QB#4	I0<3>/I0<3>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk431	I0<3>/I0<3>/I0<1>/QB#6	I0<3>/I0<3>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk432	I0<3>/I0<3>/I0<1>/QB#5	I0<3>/I0<3>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk433	I0<3>/I0<3>/I0<0>/QB#4	I0<3>/I0<3>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk434	I0<3>/I0<3>/I0<0>/QB#6	I0<3>/I0<3>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk435	I0<3>/I0<3>/I0<0>/QB#5	I0<3>/I0<3>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk436	I0<3>/I0<2>/I0<3>/QB#4	I0<3>/I0<2>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk437	I0<3>/I0<2>/I0<3>/QB#6	I0<3>/I0<2>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk438	I0<3>/I0<2>/I0<3>/QB#5	I0<3>/I0<2>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk439	I0<3>/I0<2>/I0<2>/QB#4	I0<3>/I0<2>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk440	I0<3>/I0<2>/I0<2>/QB#6	I0<3>/I0<2>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk441	I0<3>/I0<2>/I0<2>/QB#5	I0<3>/I0<2>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk442	I0<3>/I0<2>/I0<1>/QB#4	I0<3>/I0<2>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk443	I0<3>/I0<2>/I0<1>/QB#6	I0<3>/I0<2>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk444	I0<3>/I0<2>/I0<1>/QB#5	I0<3>/I0<2>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk445	I0<3>/I0<2>/I0<0>/QB#4	I0<3>/I0<2>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk446	I0<3>/I0<2>/I0<0>/QB#6	I0<3>/I0<2>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk447	I0<3>/I0<2>/I0<0>/QB#5	I0<3>/I0<2>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk448	I0<3>/I0<1>/I0<3>/QB#4	I0<3>/I0<1>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk449	I0<3>/I0<1>/I0<3>/QB#6	I0<3>/I0<1>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk450	I0<3>/I0<1>/I0<3>/QB#5	I0<3>/I0<1>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk451	I0<3>/I0<1>/I0<2>/QB#4	I0<3>/I0<1>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk452	I0<3>/I0<1>/I0<2>/QB#6	I0<3>/I0<1>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk453	I0<3>/I0<1>/I0<2>/QB#5	I0<3>/I0<1>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk454	I0<3>/I0<1>/I0<1>/QB#4	I0<3>/I0<1>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk455	I0<3>/I0<1>/I0<1>/QB#6	I0<3>/I0<1>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk456	I0<3>/I0<1>/I0<1>/QB#5	I0<3>/I0<1>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk457	I0<3>/I0<1>/I0<0>/QB#4	I0<3>/I0<1>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk458	I0<3>/I0<1>/I0<0>/QB#6	I0<3>/I0<1>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk459	I0<3>/I0<1>/I0<0>/QB#5	I0<3>/I0<1>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk460	I0<3>/I0<0>/I0<3>/QB#4	I0<3>/I0<0>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk461	I0<3>/I0<0>/I0<3>/QB#6	I0<3>/I0<0>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk462	I0<3>/I0<0>/I0<3>/QB#5	I0<3>/I0<0>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk463	I0<3>/I0<0>/I0<2>/QB#4	I0<3>/I0<0>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk464	I0<3>/I0<0>/I0<2>/QB#6	I0<3>/I0<0>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk465	I0<3>/I0<0>/I0<2>/QB#5	I0<3>/I0<0>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk466	I0<3>/I0<0>/I0<1>/QB#4	I0<3>/I0<0>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk467	I0<3>/I0<0>/I0<1>/QB#6	I0<3>/I0<0>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk468	I0<3>/I0<0>/I0<1>/QB#5	I0<3>/I0<0>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk469	I0<3>/I0<0>/I0<0>/QB#4	I0<3>/I0<0>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk470	I0<3>/I0<0>/I0<0>/QB#6	I0<3>/I0<0>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk471	I0<3>/I0<0>/I0<0>/QB#5	I0<3>/I0<0>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk472	I0<2>/I0<3>/I0<3>/QB#4	I0<2>/I0<3>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk473	I0<2>/I0<3>/I0<3>/QB#6	I0<2>/I0<3>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk474	I0<2>/I0<3>/I0<3>/QB#5	I0<2>/I0<3>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk475	I0<2>/I0<3>/I0<2>/QB#4	I0<2>/I0<3>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk476	I0<2>/I0<3>/I0<2>/QB#6	I0<2>/I0<3>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk477	I0<2>/I0<3>/I0<2>/QB#5	I0<2>/I0<3>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk478	I0<2>/I0<3>/I0<1>/QB#4	I0<2>/I0<3>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk479	I0<2>/I0<3>/I0<1>/QB#6	I0<2>/I0<3>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk480	I0<2>/I0<3>/I0<1>/QB#5	I0<2>/I0<3>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk481	I0<2>/I0<3>/I0<0>/QB#4	I0<2>/I0<3>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk482	I0<2>/I0<3>/I0<0>/QB#6	I0<2>/I0<3>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk483	I0<2>/I0<3>/I0<0>/QB#5	I0<2>/I0<3>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk484	I0<2>/I0<2>/I0<3>/QB#4	I0<2>/I0<2>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk485	I0<2>/I0<2>/I0<3>/QB#6	I0<2>/I0<2>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk486	I0<2>/I0<2>/I0<3>/QB#5	I0<2>/I0<2>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk487	I0<2>/I0<2>/I0<2>/QB#4	I0<2>/I0<2>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk488	I0<2>/I0<2>/I0<2>/QB#6	I0<2>/I0<2>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk489	I0<2>/I0<2>/I0<2>/QB#5	I0<2>/I0<2>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk490	I0<2>/I0<2>/I0<1>/QB#4	I0<2>/I0<2>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk491	I0<2>/I0<2>/I0<1>/QB#6	I0<2>/I0<2>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk492	I0<2>/I0<2>/I0<1>/QB#5	I0<2>/I0<2>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk493	I0<2>/I0<2>/I0<0>/QB#4	I0<2>/I0<2>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk494	I0<2>/I0<2>/I0<0>/QB#6	I0<2>/I0<2>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk495	I0<2>/I0<2>/I0<0>/QB#5	I0<2>/I0<2>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk496	I0<2>/I0<1>/I0<3>/QB#4	I0<2>/I0<1>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk497	I0<2>/I0<1>/I0<3>/QB#6	I0<2>/I0<1>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk498	I0<2>/I0<1>/I0<3>/QB#5	I0<2>/I0<1>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk499	I0<2>/I0<1>/I0<2>/QB#4	I0<2>/I0<1>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk500	I0<2>/I0<1>/I0<2>/QB#6	I0<2>/I0<1>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk501	I0<2>/I0<1>/I0<2>/QB#5	I0<2>/I0<1>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk502	I0<2>/I0<1>/I0<1>/QB#4	I0<2>/I0<1>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk503	I0<2>/I0<1>/I0<1>/QB#6	I0<2>/I0<1>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk504	I0<2>/I0<1>/I0<1>/QB#5	I0<2>/I0<1>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk505	I0<2>/I0<1>/I0<0>/QB#4	I0<2>/I0<1>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk506	I0<2>/I0<1>/I0<0>/QB#6	I0<2>/I0<1>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk507	I0<2>/I0<1>/I0<0>/QB#5	I0<2>/I0<1>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk508	I0<2>/I0<0>/I0<3>/QB#4	I0<2>/I0<0>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk509	I0<2>/I0<0>/I0<3>/QB#6	I0<2>/I0<0>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk510	I0<2>/I0<0>/I0<3>/QB#5	I0<2>/I0<0>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk511	I0<2>/I0<0>/I0<2>/QB#4	I0<2>/I0<0>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk512	I0<2>/I0<0>/I0<2>/QB#6	I0<2>/I0<0>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk513	I0<2>/I0<0>/I0<2>/QB#5	I0<2>/I0<0>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk514	I0<2>/I0<0>/I0<1>/QB#4	I0<2>/I0<0>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk515	I0<2>/I0<0>/I0<1>/QB#6	I0<2>/I0<0>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk516	I0<2>/I0<0>/I0<1>/QB#5	I0<2>/I0<0>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk517	I0<2>/I0<0>/I0<0>/QB#4	I0<2>/I0<0>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk518	I0<2>/I0<0>/I0<0>/QB#6	I0<2>/I0<0>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk519	I0<2>/I0<0>/I0<0>/QB#5	I0<2>/I0<0>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk520	I0<1>/I0<3>/I0<3>/QB#4	I0<1>/I0<3>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk521	I0<1>/I0<3>/I0<3>/QB#6	I0<1>/I0<3>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk522	I0<1>/I0<3>/I0<3>/QB#5	I0<1>/I0<3>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk523	I0<1>/I0<3>/I0<2>/QB#4	I0<1>/I0<3>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk524	I0<1>/I0<3>/I0<2>/QB#6	I0<1>/I0<3>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk525	I0<1>/I0<3>/I0<2>/QB#5	I0<1>/I0<3>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk526	I0<1>/I0<3>/I0<1>/QB#4	I0<1>/I0<3>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk527	I0<1>/I0<3>/I0<1>/QB#6	I0<1>/I0<3>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk528	I0<1>/I0<3>/I0<1>/QB#5	I0<1>/I0<3>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk529	I0<1>/I0<3>/I0<0>/QB#4	I0<1>/I0<3>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk530	I0<1>/I0<3>/I0<0>/QB#6	I0<1>/I0<3>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk531	I0<1>/I0<3>/I0<0>/QB#5	I0<1>/I0<3>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk532	I0<1>/I0<2>/I0<3>/QB#4	I0<1>/I0<2>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk533	I0<1>/I0<2>/I0<3>/QB#6	I0<1>/I0<2>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk534	I0<1>/I0<2>/I0<3>/QB#5	I0<1>/I0<2>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk535	I0<1>/I0<2>/I0<2>/QB#4	I0<1>/I0<2>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk536	I0<1>/I0<2>/I0<2>/QB#6	I0<1>/I0<2>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk537	I0<1>/I0<2>/I0<2>/QB#5	I0<1>/I0<2>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk538	I0<1>/I0<2>/I0<1>/QB#4	I0<1>/I0<2>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk539	I0<1>/I0<2>/I0<1>/QB#6	I0<1>/I0<2>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk540	I0<1>/I0<2>/I0<1>/QB#5	I0<1>/I0<2>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk541	I0<1>/I0<2>/I0<0>/QB#4	I0<1>/I0<2>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk542	I0<1>/I0<2>/I0<0>/QB#6	I0<1>/I0<2>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk543	I0<1>/I0<2>/I0<0>/QB#5	I0<1>/I0<2>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk544	I0<1>/I0<1>/I0<3>/QB#4	I0<1>/I0<1>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk545	I0<1>/I0<1>/I0<3>/QB#6	I0<1>/I0<1>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk546	I0<1>/I0<1>/I0<3>/QB#5	I0<1>/I0<1>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk547	I0<1>/I0<1>/I0<2>/QB#4	I0<1>/I0<1>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk548	I0<1>/I0<1>/I0<2>/QB#6	I0<1>/I0<1>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk549	I0<1>/I0<1>/I0<2>/QB#5	I0<1>/I0<1>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk550	I0<1>/I0<1>/I0<1>/QB#4	I0<1>/I0<1>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk551	I0<1>/I0<1>/I0<1>/QB#6	I0<1>/I0<1>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk552	I0<1>/I0<1>/I0<1>/QB#5	I0<1>/I0<1>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk553	I0<1>/I0<1>/I0<0>/QB#4	I0<1>/I0<1>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk554	I0<1>/I0<1>/I0<0>/QB#6	I0<1>/I0<1>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk555	I0<1>/I0<1>/I0<0>/QB#5	I0<1>/I0<1>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk556	I0<1>/I0<0>/I0<3>/QB#4	I0<1>/I0<0>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk557	I0<1>/I0<0>/I0<3>/QB#6	I0<1>/I0<0>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk558	I0<1>/I0<0>/I0<3>/QB#5	I0<1>/I0<0>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk559	I0<1>/I0<0>/I0<2>/QB#4	I0<1>/I0<0>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk560	I0<1>/I0<0>/I0<2>/QB#6	I0<1>/I0<0>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk561	I0<1>/I0<0>/I0<2>/QB#5	I0<1>/I0<0>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk562	I0<1>/I0<0>/I0<1>/QB#4	I0<1>/I0<0>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk563	I0<1>/I0<0>/I0<1>/QB#6	I0<1>/I0<0>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk564	I0<1>/I0<0>/I0<1>/QB#5	I0<1>/I0<0>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk565	I0<1>/I0<0>/I0<0>/QB#4	I0<1>/I0<0>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk566	I0<1>/I0<0>/I0<0>/QB#6	I0<1>/I0<0>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk567	I0<1>/I0<0>/I0<0>/QB#5	I0<1>/I0<0>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk568	I0<0>/I0<3>/I0<3>/QB#4	I0<0>/I0<3>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk569	I0<0>/I0<3>/I0<3>/QB#6	I0<0>/I0<3>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk570	I0<0>/I0<3>/I0<3>/QB#5	I0<0>/I0<3>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk571	I0<0>/I0<3>/I0<2>/QB#4	I0<0>/I0<3>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk572	I0<0>/I0<3>/I0<2>/QB#6	I0<0>/I0<3>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk573	I0<0>/I0<3>/I0<2>/QB#5	I0<0>/I0<3>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk574	I0<0>/I0<3>/I0<1>/QB#4	I0<0>/I0<3>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk575	I0<0>/I0<3>/I0<1>/QB#6	I0<0>/I0<3>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk576	I0<0>/I0<3>/I0<1>/QB#5	I0<0>/I0<3>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk577	I0<0>/I0<3>/I0<0>/QB#4	I0<0>/I0<3>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk578	I0<0>/I0<3>/I0<0>/QB#6	I0<0>/I0<3>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk579	I0<0>/I0<3>/I0<0>/QB#5	I0<0>/I0<3>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk580	I0<0>/I0<2>/I0<3>/QB#4	I0<0>/I0<2>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk581	I0<0>/I0<2>/I0<3>/QB#6	I0<0>/I0<2>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk582	I0<0>/I0<2>/I0<3>/QB#5	I0<0>/I0<2>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk583	I0<0>/I0<2>/I0<2>/QB#4	I0<0>/I0<2>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk584	I0<0>/I0<2>/I0<2>/QB#6	I0<0>/I0<2>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk585	I0<0>/I0<2>/I0<2>/QB#5	I0<0>/I0<2>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk586	I0<0>/I0<2>/I0<1>/QB#4	I0<0>/I0<2>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk587	I0<0>/I0<2>/I0<1>/QB#6	I0<0>/I0<2>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk588	I0<0>/I0<2>/I0<1>/QB#5	I0<0>/I0<2>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk589	I0<0>/I0<2>/I0<0>/QB#4	I0<0>/I0<2>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk590	I0<0>/I0<2>/I0<0>/QB#6	I0<0>/I0<2>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk591	I0<0>/I0<2>/I0<0>/QB#5	I0<0>/I0<2>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk592	I0<0>/I0<1>/I0<3>/QB#4	I0<0>/I0<1>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk593	I0<0>/I0<1>/I0<3>/QB#6	I0<0>/I0<1>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk594	I0<0>/I0<1>/I0<3>/QB#5	I0<0>/I0<1>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk595	I0<0>/I0<1>/I0<2>/QB#4	I0<0>/I0<1>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk596	I0<0>/I0<1>/I0<2>/QB#6	I0<0>/I0<1>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk597	I0<0>/I0<1>/I0<2>/QB#5	I0<0>/I0<1>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk598	I0<0>/I0<1>/I0<1>/QB#4	I0<0>/I0<1>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk599	I0<0>/I0<1>/I0<1>/QB#6	I0<0>/I0<1>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk600	I0<0>/I0<1>/I0<1>/QB#5	I0<0>/I0<1>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk601	I0<0>/I0<1>/I0<0>/QB#4	I0<0>/I0<1>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk602	I0<0>/I0<1>/I0<0>/QB#6	I0<0>/I0<1>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk603	I0<0>/I0<1>/I0<0>/QB#5	I0<0>/I0<1>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk604	I0<0>/I0<0>/I0<3>/QB#4	I0<0>/I0<0>/I0<3>/QB#6	   75.2879
+ $metal1_conn
Rk605	I0<0>/I0<0>/I0<3>/QB#6	I0<0>/I0<0>/I0<3>/QB	    0.1682
+ $metal1_conn
Rk606	I0<0>/I0<0>/I0<3>/QB#5	I0<0>/I0<0>/I0<3>/QB#6	   62.0000
+ $metal1_conn
Rk607	I0<0>/I0<0>/I0<2>/QB#4	I0<0>/I0<0>/I0<2>/QB#6	   75.2879
+ $metal1_conn
Rk608	I0<0>/I0<0>/I0<2>/QB#6	I0<0>/I0<0>/I0<2>/QB#3	    0.1682
+ $metal1_conn
Rk609	I0<0>/I0<0>/I0<2>/QB#5	I0<0>/I0<0>/I0<2>/QB#6	   62.0000
+ $metal1_conn
Rk610	I0<0>/I0<0>/I0<1>/QB#4	I0<0>/I0<0>/I0<1>/QB#6	   75.2879
+ $metal1_conn
Rk611	I0<0>/I0<0>/I0<1>/QB#6	I0<0>/I0<0>/I0<1>/QB	    0.1682
+ $metal1_conn
Rk612	I0<0>/I0<0>/I0<1>/QB#5	I0<0>/I0<0>/I0<1>/QB#6	   62.0000
+ $metal1_conn
Rk613	I0<0>/I0<0>/I0<0>/QB#4	I0<0>/I0<0>/I0<0>/QB#6	   75.2879
+ $metal1_conn
Rk614	I0<0>/I0<0>/I0<0>/QB#6	I0<0>/I0<0>/I0<0>/QB#3	    0.1682
+ $metal1_conn
Rk615	I0<0>/I0<0>/I0<0>/QB#5	I0<0>/I0<0>/I0<0>/QB#6	   62.0000
+ $metal1_conn
Rk616	VSS#70	VSS#1	   27.3724	$metal1_conn
Rk617	WL<63>#4	WL<63>#6	    6.6000	$metal1_conn
Rk618	WL<62>#3	WL<62>#6	    6.6000	$metal1_conn
Rk619	WL<61>#4	WL<61>#6	    6.6000	$metal1_conn
Rk620	WL<60>#3	WL<60>#6	    6.6000	$metal1_conn
Rk621	WL<59>#4	WL<59>#6	    6.6000	$metal1_conn
Rk622	WL<58>#3	WL<58>#6	    6.6000	$metal1_conn
Rk623	WL<57>#4	WL<57>#6	    6.6000	$metal1_conn
Rk624	WL<56>#3	WL<56>#6	    6.6000	$metal1_conn
Rk625	WL<55>#4	WL<55>#6	    6.6000	$metal1_conn
Rk626	WL<54>#3	WL<54>#6	    6.6000	$metal1_conn
Rk627	WL<53>#4	WL<53>#6	    6.6000	$metal1_conn
Rk628	WL<52>#3	WL<52>#6	    6.6000	$metal1_conn
Rk629	WL<51>#4	WL<51>#6	    6.6000	$metal1_conn
Rk630	WL<50>#3	WL<50>#6	    6.6000	$metal1_conn
Rk631	WL<49>#4	WL<49>#6	    6.6000	$metal1_conn
Rk632	WL<48>#3	WL<48>#6	    6.6000	$metal1_conn
Rk633	WL<47>#4	WL<47>#6	    6.6000	$metal1_conn
Rk634	WL<46>#3	WL<46>#6	    6.6000	$metal1_conn
Rk635	WL<45>#4	WL<45>#6	    6.6000	$metal1_conn
Rk636	WL<44>#3	WL<44>#6	    6.6000	$metal1_conn
Rk637	WL<43>#4	WL<43>#6	    6.6000	$metal1_conn
Rk638	WL<42>#3	WL<42>#6	    6.6000	$metal1_conn
Rk639	WL<41>#4	WL<41>#6	    6.6000	$metal1_conn
Rk640	WL<40>#3	WL<40>#6	    6.6000	$metal1_conn
Rk641	WL<39>#4	WL<39>#6	    6.6000	$metal1_conn
Rk642	WL<38>#3	WL<38>#6	    6.6000	$metal1_conn
Rk643	WL<37>#4	WL<37>#6	    6.6000	$metal1_conn
Rk644	WL<36>#3	WL<36>#6	    6.6000	$metal1_conn
Rk645	WL<35>#4	WL<35>#6	    6.6000	$metal1_conn
Rk646	WL<34>#3	WL<34>#6	    6.6000	$metal1_conn
Rk647	WL<33>#4	WL<33>#6	    6.6000	$metal1_conn
Rk648	WL<32>#3	WL<32>#6	    6.6000	$metal1_conn
Rk649	WL<31>#4	WL<31>#6	    6.6000	$metal1_conn
Rk650	WL<30>#3	WL<30>#6	    6.6000	$metal1_conn
Rk651	WL<29>#4	WL<29>#6	    6.6000	$metal1_conn
Rk652	WL<28>#3	WL<28>#6	    6.6000	$metal1_conn
Rk653	WL<27>#4	WL<27>#6	    6.6000	$metal1_conn
Rk654	WL<26>#3	WL<26>#6	    6.6000	$metal1_conn
Rk655	WL<25>#4	WL<25>#6	    6.6000	$metal1_conn
Rk656	WL<24>#3	WL<24>#6	    6.6000	$metal1_conn
Rk657	WL<23>#4	WL<23>#6	    6.6000	$metal1_conn
Rk658	WL<22>#3	WL<22>#6	    6.6000	$metal1_conn
Rk659	WL<21>#4	WL<21>#6	    6.6000	$metal1_conn
Rk660	WL<20>#3	WL<20>#6	    6.6000	$metal1_conn
Rk661	WL<19>#4	WL<19>#6	    6.6000	$metal1_conn
Rk662	WL<18>#3	WL<18>#6	    6.6000	$metal1_conn
Rk663	WL<17>#4	WL<17>#6	    6.6000	$metal1_conn
Rk664	WL<16>#3	WL<16>#6	    6.6000	$metal1_conn
Rk665	WL<15>#4	WL<15>#6	    6.6000	$metal1_conn
Rk666	WL<14>#3	WL<14>#6	    6.6000	$metal1_conn
Rk667	WL<13>#4	WL<13>#6	    6.6000	$metal1_conn
Rk668	WL<12>#3	WL<12>#6	    6.6000	$metal1_conn
Rk669	WL<11>#4	WL<11>#6	    6.6000	$metal1_conn
Rk670	WL<10>#3	WL<10>#6	    6.6000	$metal1_conn
Rk671	WL<9>#4	WL<9>#6	    6.6000	$metal1_conn
Rk672	WL<8>#3	WL<8>#6	    6.6000	$metal1_conn
Rk673	WL<7>#4	WL<7>#6	    6.6000	$metal1_conn
Rk674	WL<6>#3	WL<6>#6	    6.6000	$metal1_conn
Rk675	WL<5>#4	WL<5>#6	    6.6000	$metal1_conn
Rk676	WL<4>#3	WL<4>#6	    6.6000	$metal1_conn
Rk677	WL<3>#4	WL<3>#6	    6.6000	$metal1_conn
Rk678	WL<2>#3	WL<2>#6	    6.6000	$metal1_conn
Rk679	WL<1>#4	WL<1>#6	    6.6000	$metal1_conn
Rk680	WL<0>#3	WL<0>#6	    6.6000	$metal1_conn
Rk681	VSS#71	VSS#1	   27.3724	$metal1_conn
Rk682	VSS#72	VSS#73	   81.7666	$metal1_conn
Rk683	VSS#74	VSS#75	   81.7666	$metal1_conn
Rk684	VSS#76	VSS#77	   81.7666	$metal1_conn
Rk685	VSS#78	VSS#79	   81.7666	$metal1_conn
Rk686	VSS#80	VSS#81	   81.7666	$metal1_conn
Rk687	VSS#82	VSS#83	   81.7666	$metal1_conn
Rk688	VSS#84	VSS#85	   81.7666	$metal1_conn
Rk689	VSS#86	VSS#87	   81.7666	$metal1_conn
Rk690	VSS#88	VSS#89	   81.7666	$metal1_conn
Rk691	VSS#90	VSS#91	   81.7666	$metal1_conn
Rk692	VSS#92	VSS#93	   81.7666	$metal1_conn
Rk693	VSS#94	VSS#95	   81.7666	$metal1_conn
Rk694	VSS#96	VSS#97	   81.7666	$metal1_conn
Rk695	VSS#98	VSS#99	   81.7666	$metal1_conn
Rk696	VSS#100	VSS#101	   81.7666	$metal1_conn
Rk697	VSS#102	VSS#103	   81.7666	$metal1_conn
Rk698	VSS#104	VSS#105	   81.7666	$metal1_conn
Rk699	VSS#106	VSS#107	   81.7666	$metal1_conn
Rk700	VSS#108	VSS#109	   81.7666	$metal1_conn
Rk701	VSS#110	VSS#111	   81.7666	$metal1_conn
Rk702	VSS#112	VSS#113	   81.7666	$metal1_conn
Rk703	VSS#114	VSS#115	   81.7666	$metal1_conn
Rk704	VSS#116	VSS#117	   81.7666	$metal1_conn
Rk705	VSS#118	VSS#119	   81.7666	$metal1_conn
Rk706	VSS#120	VSS#121	   81.7666	$metal1_conn
Rk707	VSS#122	VSS#123	   81.7666	$metal1_conn
Rk708	VSS#124	VSS#125	   81.7666	$metal1_conn
Rk709	VSS#126	VSS#127	   81.7666	$metal1_conn
Rk710	VSS#128	VSS#129	   81.7666	$metal1_conn
Rk711	VSS#130	VSS#131	   81.7666	$metal1_conn
Rk712	VSS#132	VSS#133	   81.7666	$metal1_conn
Rk713	VSS#134	VSS#135	   81.7666	$metal1_conn
Rj1	VSS#5	VSS#136	    6.6000	$metal2_conn
Rj2	VSS#7	VSS#137	    6.6000	$metal2_conn
Rj3	VSS#9	VSS#138	    6.6000	$metal2_conn
Rj4	VSS#11	VSS#139	    6.6000	$metal2_conn
Rj5	VSS#13	VSS#140	    6.6000	$metal2_conn
Rj6	VSS#15	VSS#141	    6.6000	$metal2_conn
Rj7	VSS#17	VSS#142	    6.6000	$metal2_conn
Rj8	VSS#19	VSS#143	    6.6000	$metal2_conn
Rj9	VSS#21	VSS#144	    6.6000	$metal2_conn
Rj10	VSS#23	VSS#145	    6.6000	$metal2_conn
Rj11	VSS#25	VSS#146	    6.6000	$metal2_conn
Rj12	VSS#27	VSS#147	    6.6000	$metal2_conn
Rj13	VSS#29	VSS#148	    6.6000	$metal2_conn
Rj14	VSS#31	VSS#149	    6.6000	$metal2_conn
Rj15	VSS#33	VSS#150	    6.6000	$metal2_conn
Rj16	VSS#35	VSS#151	    6.6000	$metal2_conn
Rj17	VSS#37	VSS#152	    6.6000	$metal2_conn
Rj18	VSS#39	VSS#153	    6.6000	$metal2_conn
Rj19	VSS#41	VSS#154	    6.6000	$metal2_conn
Rj20	VSS#43	VSS#155	    6.6000	$metal2_conn
Rj21	VSS#45	VSS#156	    6.6000	$metal2_conn
Rj22	VSS#47	VSS#157	    6.6000	$metal2_conn
Rj23	VSS#49	VSS#158	    6.6000	$metal2_conn
Rj24	VSS#51	VSS#159	    6.6000	$metal2_conn
Rj25	VSS#53	VSS#160	    6.6000	$metal2_conn
Rj26	VSS#55	VSS#161	    6.6000	$metal2_conn
Rj27	VSS#57	VSS#162	    6.6000	$metal2_conn
Rj28	VSS#59	VSS#163	    6.6000	$metal2_conn
Rj29	VSS#61	VSS#164	    6.6000	$metal2_conn
Rj30	VSS#63	VSS#165	    6.6000	$metal2_conn
Rj31	VSS#65	VSS#166	    6.6000	$metal2_conn
Rj32	VSS#67	VSS#167	    6.6000	$metal2_conn
Rj33	VSS#168	VSS#69	    6.6000	$metal2_conn
Rj34	BL#65	BL#2	    6.6000	$metal2_conn
Rj35	BL#4	BL#66	    6.6000	$metal2_conn
Rj36	BL#67	BL#6	    6.6000	$metal2_conn
Rj37	BL#8	BL#68	    6.6000	$metal2_conn
Rj38	BL#69	BL#10	    6.6000	$metal2_conn
Rj39	BL#12	BL#70	    6.6000	$metal2_conn
Rj40	BL#71	BL#14	    6.6000	$metal2_conn
Rj41	BL#16	BL#72	    6.6000	$metal2_conn
Rj42	BL#73	BL#18	    6.6000	$metal2_conn
Rj43	BL#20	BL#74	    6.6000	$metal2_conn
Rj44	BL#75	BL#22	    6.6000	$metal2_conn
Rj45	BL#24	BL#76	    6.6000	$metal2_conn
Rj46	BL#77	BL#26	    6.6000	$metal2_conn
Rj47	BL#28	BL#78	    6.6000	$metal2_conn
Rj48	BL#79	BL#30	    6.6000	$metal2_conn
Rj49	BL#32	BL#80	    6.6000	$metal2_conn
Rj50	BL#81	BL#34	    6.6000	$metal2_conn
Rj51	BL#36	BL#82	    6.6000	$metal2_conn
Rj52	BL#83	BL#38	    6.6000	$metal2_conn
Rj53	BL#40	BL#84	    6.6000	$metal2_conn
Rj54	BL#85	BL#42	    6.6000	$metal2_conn
Rj55	BL#44	BL#86	    6.6000	$metal2_conn
Rj56	BL#87	BL#46	    6.6000	$metal2_conn
Rj57	BL#48	BL#88	    6.6000	$metal2_conn
Rj58	BL#89	BL#50	    6.6000	$metal2_conn
Rj59	BL#52	BL#90	    6.6000	$metal2_conn
Rj60	BL#91	BL#54	    6.6000	$metal2_conn
Rj61	BL#56	BL#92	    6.6000	$metal2_conn
Rj62	BL#93	BL#58	    6.6000	$metal2_conn
Rj63	BL#60	BL#94	    6.6000	$metal2_conn
Rj64	BL#95	BL#62	    6.6000	$metal2_conn
Rj65	BL#64	BL#96	    6.6000	$metal2_conn
Rj66	VDD#134	VDD#1	    6.6000	$metal2_conn
Rj67	VDD#71	VDD#135	    6.6000	$metal2_conn
Rj68	VDD#136	VDD#3	    6.6000	$metal2_conn
Rj69	VDD#73	VDD#137	    6.6000	$metal2_conn
Rj70	VDD#138	VDD#5	    6.6000	$metal2_conn
Rj71	VDD#75	VDD#139	    6.6000	$metal2_conn
Rj72	VDD#140	VDD#7	    6.6000	$metal2_conn
Rj73	VDD#77	VDD#141	    6.6000	$metal2_conn
Rj74	VDD#142	VDD#9	    6.6000	$metal2_conn
Rj75	VDD#79	VDD#143	    6.6000	$metal2_conn
Rj76	VDD#144	VDD#11	    6.6000	$metal2_conn
Rj77	VDD#81	VDD#145	    6.6000	$metal2_conn
Rj78	VDD#146	VDD#13	    6.6000	$metal2_conn
Rj79	VDD#83	VDD#147	    6.6000	$metal2_conn
Rj80	VDD#148	VDD#15	    6.6000	$metal2_conn
Rj81	VDD#85	VDD#149	    6.6000	$metal2_conn
Rj82	VDD#150	VDD#17	    6.6000	$metal2_conn
Rj83	VDD#87	VDD#151	    6.6000	$metal2_conn
Rj84	VDD#152	VDD#19	    6.6000	$metal2_conn
Rj85	VDD#89	VDD#153	    6.6000	$metal2_conn
Rj86	VDD#154	VDD#21	    6.6000	$metal2_conn
Rj87	VDD#91	VDD#155	    6.6000	$metal2_conn
Rj88	VDD#156	VDD#23	    6.6000	$metal2_conn
Rj89	VDD#93	VDD#157	    6.6000	$metal2_conn
Rj90	VDD#158	VDD#25	    6.6000	$metal2_conn
Rj91	VDD#95	VDD#159	    6.6000	$metal2_conn
Rj92	VDD#160	VDD#27	    6.6000	$metal2_conn
Rj93	VDD#97	VDD#161	    6.6000	$metal2_conn
Rj94	VDD#162	VDD#29	    6.6000	$metal2_conn
Rj95	VDD#99	VDD#163	    6.6000	$metal2_conn
Rj96	VDD#164	VDD#31	    6.6000	$metal2_conn
Rj97	VDD#101	VDD#165	    6.6000	$metal2_conn
Rj98	VDD#166	VDD#33	    6.6000	$metal2_conn
Rj99	VDD#103	VDD#167	    6.6000	$metal2_conn
Rj100	VDD#168	VDD#35	    6.6000	$metal2_conn
Rj101	VDD#105	VDD#169	    6.6000	$metal2_conn
Rj102	VDD#170	VDD#37	    6.6000	$metal2_conn
Rj103	VDD#107	VDD#171	    6.6000	$metal2_conn
Rj104	VDD#172	VDD#39	    6.6000	$metal2_conn
Rj105	VDD#109	VDD#173	    6.6000	$metal2_conn
Rj106	VDD#174	VDD#41	    6.6000	$metal2_conn
Rj107	VDD#111	VDD#175	    6.6000	$metal2_conn
Rj108	VDD#176	VDD#43	    6.6000	$metal2_conn
Rj109	VDD#113	VDD#177	    6.6000	$metal2_conn
Rj110	VDD#178	VDD#45	    6.6000	$metal2_conn
Rj111	VDD#115	VDD#179	    6.6000	$metal2_conn
Rj112	VDD#180	VDD#47	    6.6000	$metal2_conn
Rj113	VDD#117	VDD#181	    6.6000	$metal2_conn
Rj114	VDD#182	VDD#49	    6.6000	$metal2_conn
Rj115	VDD#119	VDD#183	    6.6000	$metal2_conn
Rj116	VDD#184	VDD#51	    6.6000	$metal2_conn
Rj117	VDD#121	VDD#185	    6.6000	$metal2_conn
Rj118	VDD#186	VDD#53	    6.6000	$metal2_conn
Rj119	VDD#123	VDD#187	    6.6000	$metal2_conn
Rj120	VDD#188	VDD#55	    6.6000	$metal2_conn
Rj121	VDD#125	VDD#189	    6.6000	$metal2_conn
Rj122	VDD#190	VDD#57	    6.6000	$metal2_conn
Rj123	VDD#127	VDD#191	    6.6000	$metal2_conn
Rj124	VDD#192	VDD#59	    6.6000	$metal2_conn
Rj125	VDD#129	VDD#193	    6.6000	$metal2_conn
Rj126	VDD#194	VDD#61	    6.6000	$metal2_conn
Rj127	VDD#131	VDD#195	    6.6000	$metal2_conn
Rj128	VDD#196	VDD#63	    6.6000	$metal2_conn
Rj129	VDD#133	VDD#197	    6.6000	$metal2_conn
Rj130	VDD#198	VDD#65	    6.6000	$metal2_conn
Rj131	BLB#67	BLB#2	    6.6000	$metal2_conn
Rj132	BLB#4	BLB#68	    6.6000	$metal2_conn
Rj133	BLB#69	BLB#6	    6.6000	$metal2_conn
Rj134	BLB#8	BLB#70	    6.6000	$metal2_conn
Rj135	BLB#71	BLB#10	    6.6000	$metal2_conn
Rj136	BLB#12	BLB#72	    6.6000	$metal2_conn
Rj137	BLB#73	BLB#14	    6.6000	$metal2_conn
Rj138	BLB#16	BLB#74	    6.6000	$metal2_conn
Rj139	BLB#75	BLB#18	    6.6000	$metal2_conn
Rj140	BLB#20	BLB#76	    6.6000	$metal2_conn
Rj141	BLB#77	BLB#22	    6.6000	$metal2_conn
Rj142	BLB#24	BLB#78	    6.6000	$metal2_conn
Rj143	BLB#79	BLB#26	    6.6000	$metal2_conn
Rj144	BLB#28	BLB#80	    6.6000	$metal2_conn
Rj145	BLB#81	BLB#30	    6.6000	$metal2_conn
Rj146	BLB#32	BLB#82	    6.6000	$metal2_conn
Rj147	BLB#83	BLB#34	    6.6000	$metal2_conn
Rj148	BLB#36	BLB#84	    6.6000	$metal2_conn
Rj149	BLB#85	BLB#38	    6.6000	$metal2_conn
Rj150	BLB#40	BLB#86	    6.6000	$metal2_conn
Rj151	BLB#87	BLB#42	    6.6000	$metal2_conn
Rj152	BLB#44	BLB#88	    6.6000	$metal2_conn
Rj153	BLB#89	BLB#46	    6.6000	$metal2_conn
Rj154	BLB#48	BLB#90	    6.6000	$metal2_conn
Rj155	BLB#91	BLB#50	    6.6000	$metal2_conn
Rj156	BLB#52	BLB#92	    6.6000	$metal2_conn
Rj157	BLB#93	BLB#54	    6.6000	$metal2_conn
Rj158	BLB#56	BLB#94	    6.6000	$metal2_conn
Rj159	BLB#95	BLB#58	    6.6000	$metal2_conn
Rj160	BLB#60	BLB#96	    6.6000	$metal2_conn
Rj161	BLB#97	BLB#62	    6.6000	$metal2_conn
Rj162	BLB#64	BLB#98	    6.6000	$metal2_conn
Rj163	BLB#99	BLB#66	    6.6000	$metal2_conn
Rj164	VDD#67	VDD#199	    6.6000	$metal2_conn
Rj165	VDD#69	VDD#200	    6.6000	$metal2_conn
Rj167	VSS#70	VSS#2	    0.9767	$metal2_conn
Rj168	VSS#2	VSS#170	    6.6000	$metal2_conn
Rj170	VSS#71	VSS#3	    0.9767	$metal2_conn
Rj172	WL<63>#6	WL<63>#7	    0.9163	$metal2_conn
Rj173	WL<63>#7	WL<63>	4.614e-02	$metal2_conn
Rj174	WL<63>#7	WL<63>#5	3.578e-02	$metal2_conn
Rj175	WL<62>#6	WL<62>#7	    0.9163	$metal2_conn
Rj176	WL<62>#7	WL<62>	4.614e-02	$metal2_conn
Rj177	WL<62>#7	WL<62>#5	3.578e-02	$metal2_conn
Rj178	WL<61>#6	WL<61>#7	    0.9163	$metal2_conn
Rj179	WL<61>#7	WL<61>	4.614e-02	$metal2_conn
Rj180	WL<61>#7	WL<61>#5	3.578e-02	$metal2_conn
Rj181	WL<60>#6	WL<60>#7	    0.9163	$metal2_conn
Rj182	WL<60>#7	WL<60>	4.614e-02	$metal2_conn
Rj183	WL<60>#7	WL<60>#5	3.578e-02	$metal2_conn
Rj184	WL<59>#6	WL<59>#7	    0.9163	$metal2_conn
Rj185	WL<59>#7	WL<59>	4.614e-02	$metal2_conn
Rj186	WL<59>#7	WL<59>#5	3.578e-02	$metal2_conn
Rj187	WL<58>#6	WL<58>#7	    0.9163	$metal2_conn
Rj188	WL<58>#7	WL<58>	4.614e-02	$metal2_conn
Rj189	WL<58>#7	WL<58>#5	3.578e-02	$metal2_conn
Rj190	WL<57>#6	WL<57>#7	    0.9163	$metal2_conn
Rj191	WL<57>#7	WL<57>	4.614e-02	$metal2_conn
Rj192	WL<57>#7	WL<57>#5	3.578e-02	$metal2_conn
Rj193	WL<56>#6	WL<56>#7	    0.9163	$metal2_conn
Rj194	WL<56>#7	WL<56>	4.614e-02	$metal2_conn
Rj195	WL<56>#7	WL<56>#5	3.578e-02	$metal2_conn
Rj196	WL<55>#6	WL<55>#7	    0.9163	$metal2_conn
Rj197	WL<55>#7	WL<55>	4.614e-02	$metal2_conn
Rj198	WL<55>#7	WL<55>#5	3.578e-02	$metal2_conn
Rj199	WL<54>#6	WL<54>#7	    0.9163	$metal2_conn
Rj200	WL<54>#7	WL<54>	4.614e-02	$metal2_conn
Rj201	WL<54>#7	WL<54>#5	3.578e-02	$metal2_conn
Rj202	WL<53>#6	WL<53>#7	    0.9163	$metal2_conn
Rj203	WL<53>#7	WL<53>	4.614e-02	$metal2_conn
Rj204	WL<53>#7	WL<53>#5	3.578e-02	$metal2_conn
Rj205	WL<52>#6	WL<52>#7	    0.9163	$metal2_conn
Rj206	WL<52>#7	WL<52>	4.614e-02	$metal2_conn
Rj207	WL<52>#7	WL<52>#5	3.578e-02	$metal2_conn
Rj208	WL<51>#6	WL<51>#7	    0.9163	$metal2_conn
Rj209	WL<51>#7	WL<51>	4.614e-02	$metal2_conn
Rj210	WL<51>#7	WL<51>#5	3.578e-02	$metal2_conn
Rj211	WL<50>#6	WL<50>#7	    0.9163	$metal2_conn
Rj212	WL<50>#7	WL<50>	4.614e-02	$metal2_conn
Rj213	WL<50>#7	WL<50>#5	3.578e-02	$metal2_conn
Rj214	WL<49>#6	WL<49>#7	    0.9163	$metal2_conn
Rj215	WL<49>#7	WL<49>	4.614e-02	$metal2_conn
Rj216	WL<49>#7	WL<49>#5	3.578e-02	$metal2_conn
Rj217	WL<48>#6	WL<48>#7	    0.9163	$metal2_conn
Rj218	WL<48>#7	WL<48>	4.614e-02	$metal2_conn
Rj219	WL<48>#7	WL<48>#5	3.578e-02	$metal2_conn
Rj220	WL<47>#6	WL<47>#7	    0.9163	$metal2_conn
Rj221	WL<47>#7	WL<47>	4.614e-02	$metal2_conn
Rj222	WL<47>#7	WL<47>#5	3.578e-02	$metal2_conn
Rj223	WL<46>#6	WL<46>#7	    0.9163	$metal2_conn
Rj224	WL<46>#7	WL<46>	4.614e-02	$metal2_conn
Rj225	WL<46>#7	WL<46>#5	3.578e-02	$metal2_conn
Rj226	WL<45>#6	WL<45>#7	    0.9163	$metal2_conn
Rj227	WL<45>#7	WL<45>	4.614e-02	$metal2_conn
Rj228	WL<45>#7	WL<45>#5	3.578e-02	$metal2_conn
Rj229	WL<44>#6	WL<44>#7	    0.9163	$metal2_conn
Rj230	WL<44>#7	WL<44>	4.614e-02	$metal2_conn
Rj231	WL<44>#7	WL<44>#5	3.578e-02	$metal2_conn
Rj232	WL<43>#6	WL<43>#7	    0.9163	$metal2_conn
Rj233	WL<43>#7	WL<43>	4.614e-02	$metal2_conn
Rj234	WL<43>#7	WL<43>#5	3.578e-02	$metal2_conn
Rj235	WL<42>#6	WL<42>#7	    0.9163	$metal2_conn
Rj236	WL<42>#7	WL<42>	4.614e-02	$metal2_conn
Rj237	WL<42>#7	WL<42>#5	3.578e-02	$metal2_conn
Rj238	WL<41>#6	WL<41>#7	    0.9163	$metal2_conn
Rj239	WL<41>#7	WL<41>	4.614e-02	$metal2_conn
Rj240	WL<41>#7	WL<41>#5	3.578e-02	$metal2_conn
Rj241	WL<40>#6	WL<40>#7	    0.9163	$metal2_conn
Rj242	WL<40>#7	WL<40>	4.614e-02	$metal2_conn
Rj243	WL<40>#7	WL<40>#5	3.578e-02	$metal2_conn
Rj244	WL<39>#6	WL<39>#7	    0.9163	$metal2_conn
Rj245	WL<39>#7	WL<39>	4.614e-02	$metal2_conn
Rj246	WL<39>#7	WL<39>#5	3.578e-02	$metal2_conn
Rj247	WL<38>#6	WL<38>#7	    0.9163	$metal2_conn
Rj248	WL<38>#7	WL<38>	4.614e-02	$metal2_conn
Rj249	WL<38>#7	WL<38>#5	3.578e-02	$metal2_conn
Rj250	WL<37>#6	WL<37>#7	    0.9163	$metal2_conn
Rj251	WL<37>#7	WL<37>	4.614e-02	$metal2_conn
Rj252	WL<37>#7	WL<37>#5	3.578e-02	$metal2_conn
Rj253	WL<36>#6	WL<36>#7	    0.9163	$metal2_conn
Rj254	WL<36>#7	WL<36>	4.614e-02	$metal2_conn
Rj255	WL<36>#7	WL<36>#5	3.578e-02	$metal2_conn
Rj256	WL<35>#6	WL<35>#7	    0.9163	$metal2_conn
Rj257	WL<35>#7	WL<35>	4.614e-02	$metal2_conn
Rj258	WL<35>#7	WL<35>#5	3.578e-02	$metal2_conn
Rj259	WL<34>#6	WL<34>#7	    0.9163	$metal2_conn
Rj260	WL<34>#7	WL<34>	4.614e-02	$metal2_conn
Rj261	WL<34>#7	WL<34>#5	3.578e-02	$metal2_conn
Rj262	WL<33>#6	WL<33>#7	    0.9163	$metal2_conn
Rj263	WL<33>#7	WL<33>	4.614e-02	$metal2_conn
Rj264	WL<33>#7	WL<33>#5	3.578e-02	$metal2_conn
Rj265	WL<32>#6	WL<32>#7	    0.9163	$metal2_conn
Rj266	WL<32>#7	WL<32>	4.614e-02	$metal2_conn
Rj267	WL<32>#7	WL<32>#5	3.578e-02	$metal2_conn
Rj268	WL<31>#6	WL<31>#7	    0.9163	$metal2_conn
Rj269	WL<31>#7	WL<31>	4.614e-02	$metal2_conn
Rj270	WL<31>#7	WL<31>#5	3.578e-02	$metal2_conn
Rj271	WL<30>#6	WL<30>#7	    0.9163	$metal2_conn
Rj272	WL<30>#7	WL<30>	4.614e-02	$metal2_conn
Rj273	WL<30>#7	WL<30>#5	3.578e-02	$metal2_conn
Rj274	WL<29>#6	WL<29>#7	    0.9163	$metal2_conn
Rj275	WL<29>#7	WL<29>	4.614e-02	$metal2_conn
Rj276	WL<29>#7	WL<29>#5	3.578e-02	$metal2_conn
Rj277	WL<28>#6	WL<28>#7	    0.9163	$metal2_conn
Rj278	WL<28>#7	WL<28>	4.614e-02	$metal2_conn
Rj279	WL<28>#7	WL<28>#5	3.578e-02	$metal2_conn
Rj280	WL<27>#6	WL<27>#7	    0.9163	$metal2_conn
Rj281	WL<27>#7	WL<27>	4.614e-02	$metal2_conn
Rj282	WL<27>#7	WL<27>#5	3.578e-02	$metal2_conn
Rj283	WL<26>#6	WL<26>#7	    0.9163	$metal2_conn
Rj284	WL<26>#7	WL<26>	4.614e-02	$metal2_conn
Rj285	WL<26>#7	WL<26>#5	3.578e-02	$metal2_conn
Rj286	WL<25>#6	WL<25>#7	    0.9163	$metal2_conn
Rj287	WL<25>#7	WL<25>	4.614e-02	$metal2_conn
Rj288	WL<25>#7	WL<25>#5	3.578e-02	$metal2_conn
Rj289	WL<24>#6	WL<24>#7	    0.9163	$metal2_conn
Rj290	WL<24>#7	WL<24>	4.614e-02	$metal2_conn
Rj291	WL<24>#7	WL<24>#5	3.578e-02	$metal2_conn
Rj292	WL<23>#6	WL<23>#7	    0.9163	$metal2_conn
Rj293	WL<23>#7	WL<23>	4.614e-02	$metal2_conn
Rj294	WL<23>#7	WL<23>#5	3.578e-02	$metal2_conn
Rj295	WL<22>#6	WL<22>#7	    0.9163	$metal2_conn
Rj296	WL<22>#7	WL<22>	4.614e-02	$metal2_conn
Rj297	WL<22>#7	WL<22>#5	3.578e-02	$metal2_conn
Rj298	WL<21>#6	WL<21>#7	    0.9163	$metal2_conn
Rj299	WL<21>#7	WL<21>	4.614e-02	$metal2_conn
Rj300	WL<21>#7	WL<21>#5	3.578e-02	$metal2_conn
Rj301	WL<20>#6	WL<20>#7	    0.9163	$metal2_conn
Rj302	WL<20>#7	WL<20>	4.614e-02	$metal2_conn
Rj303	WL<20>#7	WL<20>#5	3.578e-02	$metal2_conn
Rj304	WL<19>#6	WL<19>#7	    0.9163	$metal2_conn
Rj305	WL<19>#7	WL<19>	4.614e-02	$metal2_conn
Rj306	WL<19>#7	WL<19>#5	3.578e-02	$metal2_conn
Rj307	WL<18>#6	WL<18>#7	    0.9163	$metal2_conn
Rj308	WL<18>#7	WL<18>	4.614e-02	$metal2_conn
Rj309	WL<18>#7	WL<18>#5	3.578e-02	$metal2_conn
Rj310	WL<17>#6	WL<17>#7	    0.9163	$metal2_conn
Rj311	WL<17>#7	WL<17>	4.614e-02	$metal2_conn
Rj312	WL<17>#7	WL<17>#5	3.578e-02	$metal2_conn
Rj313	WL<16>#6	WL<16>#7	    0.9163	$metal2_conn
Rj314	WL<16>#7	WL<16>	4.614e-02	$metal2_conn
Rj315	WL<16>#7	WL<16>#5	3.578e-02	$metal2_conn
Rj316	WL<15>#6	WL<15>#7	    0.9163	$metal2_conn
Rj317	WL<15>#7	WL<15>	4.614e-02	$metal2_conn
Rj318	WL<15>#7	WL<15>#5	3.578e-02	$metal2_conn
Rj319	WL<14>#6	WL<14>#7	    0.9163	$metal2_conn
Rj320	WL<14>#7	WL<14>	4.614e-02	$metal2_conn
Rj321	WL<14>#7	WL<14>#5	3.578e-02	$metal2_conn
Rj322	WL<13>#6	WL<13>#7	    0.9163	$metal2_conn
Rj323	WL<13>#7	WL<13>	4.614e-02	$metal2_conn
Rj324	WL<13>#7	WL<13>#5	3.578e-02	$metal2_conn
Rj325	WL<12>#6	WL<12>#7	    0.9163	$metal2_conn
Rj326	WL<12>#7	WL<12>	4.614e-02	$metal2_conn
Rj327	WL<12>#7	WL<12>#5	3.578e-02	$metal2_conn
Rj328	WL<11>#6	WL<11>#7	    0.9163	$metal2_conn
Rj329	WL<11>#7	WL<11>	4.614e-02	$metal2_conn
Rj330	WL<11>#7	WL<11>#5	3.578e-02	$metal2_conn
Rj331	WL<10>#6	WL<10>#7	    0.9163	$metal2_conn
Rj332	WL<10>#7	WL<10>	4.614e-02	$metal2_conn
Rj333	WL<10>#7	WL<10>#5	3.578e-02	$metal2_conn
Rj334	WL<9>#6	WL<9>#7	    0.9163	$metal2_conn
Rj335	WL<9>#7	WL<9>	4.614e-02	$metal2_conn
Rj336	WL<9>#7	WL<9>#5	3.578e-02	$metal2_conn
Rj337	WL<8>#6	WL<8>#7	    0.9163	$metal2_conn
Rj338	WL<8>#7	WL<8>	4.614e-02	$metal2_conn
Rj339	WL<8>#7	WL<8>#5	3.578e-02	$metal2_conn
Rj340	WL<7>#6	WL<7>#7	    0.9163	$metal2_conn
Rj341	WL<7>#7	WL<7>	4.614e-02	$metal2_conn
Rj342	WL<7>#7	WL<7>#5	3.578e-02	$metal2_conn
Rj343	WL<6>#6	WL<6>#7	    0.9163	$metal2_conn
Rj344	WL<6>#7	WL<6>	4.614e-02	$metal2_conn
Rj345	WL<6>#7	WL<6>#5	3.578e-02	$metal2_conn
Rj346	WL<5>#6	WL<5>#7	    0.9163	$metal2_conn
Rj347	WL<5>#7	WL<5>	4.614e-02	$metal2_conn
Rj348	WL<5>#7	WL<5>#5	3.578e-02	$metal2_conn
Rj349	WL<4>#6	WL<4>#7	    0.9163	$metal2_conn
Rj350	WL<4>#7	WL<4>	4.614e-02	$metal2_conn
Rj351	WL<4>#7	WL<4>#5	3.578e-02	$metal2_conn
Rj352	WL<3>#6	WL<3>#7	    0.9163	$metal2_conn
Rj353	WL<3>#7	WL<3>	4.614e-02	$metal2_conn
Rj354	WL<3>#7	WL<3>#5	3.578e-02	$metal2_conn
Rj355	WL<2>#6	WL<2>#7	    0.9163	$metal2_conn
Rj356	WL<2>#7	WL<2>	4.614e-02	$metal2_conn
Rj357	WL<2>#7	WL<2>#5	3.578e-02	$metal2_conn
Rj358	WL<1>#6	WL<1>#7	    0.9163	$metal2_conn
Rj359	WL<1>#7	WL<1>	4.614e-02	$metal2_conn
Rj360	WL<1>#7	WL<1>#5	3.578e-02	$metal2_conn
Rj361	WL<0>#6	WL<0>#7	    0.9163	$metal2_conn
Rj362	WL<0>#7	WL<0>	4.614e-02	$metal2_conn
Rj363	WL<0>#7	WL<0>#5	3.578e-02	$metal2_conn
Rj364	VSS#72	VSS#173	    6.6000	$metal2_conn
Rj365	VSS#74	VSS#174	    6.6000	$metal2_conn
Rj366	VSS#76	VSS#175	    6.6000	$metal2_conn
Rj367	VSS#78	VSS#176	    6.6000	$metal2_conn
Rj368	VSS#80	VSS#177	    6.6000	$metal2_conn
Rj369	VSS#82	VSS#178	    6.6000	$metal2_conn
Rj370	VSS#84	VSS#179	    6.6000	$metal2_conn
Rj371	VSS#86	VSS#180	    6.6000	$metal2_conn
Rj372	VSS#88	VSS#181	    6.6000	$metal2_conn
Rj373	VSS#90	VSS#182	    6.6000	$metal2_conn
Rj374	VSS#92	VSS#183	    6.6000	$metal2_conn
Rj375	VSS#94	VSS#184	    6.6000	$metal2_conn
Rj376	VSS#96	VSS#185	    6.6000	$metal2_conn
Rj377	VSS#98	VSS#186	    6.6000	$metal2_conn
Rj378	VSS#100	VSS#187	    6.6000	$metal2_conn
Rj379	VSS#102	VSS#188	    6.6000	$metal2_conn
Rj380	VSS#104	VSS#189	    6.6000	$metal2_conn
Rj381	VSS#106	VSS#190	    6.6000	$metal2_conn
Rj382	VSS#108	VSS#191	    6.6000	$metal2_conn
Rj383	VSS#110	VSS#192	    6.6000	$metal2_conn
Rj384	VSS#112	VSS#193	    6.6000	$metal2_conn
Rj385	VSS#114	VSS#194	    6.6000	$metal2_conn
Rj386	VSS#116	VSS#195	    6.6000	$metal2_conn
Rj387	VSS#118	VSS#196	    6.6000	$metal2_conn
Rj388	VSS#120	VSS#197	    6.6000	$metal2_conn
Rj389	VSS#122	VSS#198	    6.6000	$metal2_conn
Rj390	VSS#124	VSS#199	    6.6000	$metal2_conn
Rj391	VSS#126	VSS#200	    6.6000	$metal2_conn
Rj392	VSS#128	VSS#201	    6.6000	$metal2_conn
Rj393	VSS#130	VSS#202	    6.6000	$metal2_conn
Rj394	VSS#132	VSS#203	    6.6000	$metal2_conn
Rj395	VSS#134	VSS#204	    6.6000	$metal2_conn
Ri1	VSS	VSS#139	    0.3833	$metal3_conn
Ri2	VSS#139	VSS#140	    0.4228	$metal3_conn
Ri3	VSS#140	VSS#141	    0.4228	$metal3_conn
Ri4	VSS#141	VSS#142	    0.4228	$metal3_conn
Ri5	VSS#142	VSS#143	    0.4228	$metal3_conn
Ri6	VSS#143	VSS#144	    0.4228	$metal3_conn
Ri7	VSS#144	VSS#145	    0.4228	$metal3_conn
Ri8	VSS#145	VSS#146	    0.4228	$metal3_conn
Ri9	VSS#146	VSS#147	    0.4228	$metal3_conn
Ri10	VSS#147	VSS#148	    0.4228	$metal3_conn
Ri11	VSS#148	VSS#149	    0.4228	$metal3_conn
Ri12	VSS#149	VSS#150	    0.4228	$metal3_conn
Ri13	VSS#150	VSS#151	    0.4228	$metal3_conn
Ri14	VSS#151	VSS#152	    0.4228	$metal3_conn
Ri15	VSS#152	VSS#153	    0.4228	$metal3_conn
Ri16	VSS#153	VSS#154	    0.4228	$metal3_conn
Ri17	VSS#154	VSS#155	    0.4228	$metal3_conn
Ri18	VSS#155	VSS#156	    0.4228	$metal3_conn
Ri19	VSS#156	VSS#157	    0.4228	$metal3_conn
Ri20	VSS#157	VSS#158	    0.4228	$metal3_conn
Ri21	VSS#158	VSS#159	    0.4228	$metal3_conn
Ri22	VSS#159	VSS#160	    0.4228	$metal3_conn
Ri23	VSS#160	VSS#161	    0.4228	$metal3_conn
Ri24	VSS#161	VSS#162	    0.4228	$metal3_conn
Ri25	VSS#162	VSS#163	    0.4228	$metal3_conn
Ri26	VSS#163	VSS#164	    0.4228	$metal3_conn
Ri27	VSS#164	VSS#165	    0.4228	$metal3_conn
Ri28	VSS#165	VSS#166	    0.4228	$metal3_conn
Ri29	VSS#166	VSS#167	    0.4228	$metal3_conn
Ri30	VSS#167	VSS#168	    0.4228	$metal3_conn
Ri31	VSS#168	VSS#3	    6.8018	$metal3_conn
Ri32	VSS	VSS#138	3.954e-02	$metal3_conn
Ri33	VSS#138	VSS#137	    0.4228	$metal3_conn
Ri34	VSS#137	VSS#136	    0.4228	$metal3_conn
Ri35	VSS#136	VSS#170	    0.2018	$metal3_conn
Ri36	BL	BL#67	    0.1672	$metal3_conn
Ri37	BL#67	BL#68	    0.4228	$metal3_conn
Ri38	BL#68	BL#69	    0.4228	$metal3_conn
Ri39	BL#69	BL#70	    0.4228	$metal3_conn
Ri40	BL#70	BL#71	    0.4228	$metal3_conn
Ri41	BL#71	BL#72	    0.4228	$metal3_conn
Ri42	BL#72	BL#73	    0.4228	$metal3_conn
Ri43	BL#73	BL#74	    0.4228	$metal3_conn
Ri44	BL#74	BL#75	    0.4228	$metal3_conn
Ri45	BL#75	BL#76	    0.4228	$metal3_conn
Ri46	BL#76	BL#77	    0.4228	$metal3_conn
Ri47	BL#77	BL#78	    0.4228	$metal3_conn
Ri48	BL#78	BL#79	    0.4228	$metal3_conn
Ri49	BL#79	BL#80	    0.4228	$metal3_conn
Ri50	BL#80	BL#81	    0.4228	$metal3_conn
Ri51	BL#81	BL#82	    0.4228	$metal3_conn
Ri52	BL#82	BL#83	    0.4228	$metal3_conn
Ri53	BL#83	BL#84	    0.4228	$metal3_conn
Ri54	BL#84	BL#85	    0.4228	$metal3_conn
Ri55	BL#85	BL#86	    0.4228	$metal3_conn
Ri56	BL#86	BL#87	    0.4228	$metal3_conn
Ri57	BL#87	BL#88	    0.4228	$metal3_conn
Ri58	BL#88	BL#89	    0.4228	$metal3_conn
Ri59	BL#89	BL#90	    0.4228	$metal3_conn
Ri60	BL#90	BL#91	    0.4228	$metal3_conn
Ri61	BL#91	BL#92	    0.4228	$metal3_conn
Ri62	BL#92	BL#93	    0.4228	$metal3_conn
Ri63	BL#93	BL#94	    0.4228	$metal3_conn
Ri64	BL#94	BL#95	    0.4228	$metal3_conn
Ri65	BL#95	BL#96	    0.4324	$metal3_conn
Ri66	BL	BL#66	    0.2556	$metal3_conn
Ri67	BL#66	BL#65	    0.4253	$metal3_conn
Ri68	VDD	VDD#139	    0.1672	$metal3_conn
Ri69	VDD#139	VDD#140	    0.2068	$metal3_conn
Ri70	VDD#140	VDD#141	    0.2068	$metal3_conn
Ri71	VDD#141	VDD#142	    0.2068	$metal3_conn
Ri72	VDD#142	VDD#143	    0.2068	$metal3_conn
Ri73	VDD#143	VDD#144	    0.2068	$metal3_conn
Ri74	VDD#144	VDD#145	    0.2068	$metal3_conn
Ri75	VDD#145	VDD#146	    0.2068	$metal3_conn
Ri76	VDD#146	VDD#147	    0.2068	$metal3_conn
Ri77	VDD#147	VDD#148	    0.2068	$metal3_conn
Ri78	VDD#148	VDD#149	    0.2068	$metal3_conn
Ri79	VDD#149	VDD#150	    0.2068	$metal3_conn
Ri80	VDD#150	VDD#151	    0.2068	$metal3_conn
Ri81	VDD#151	VDD#152	    0.2068	$metal3_conn
Ri82	VDD#152	VDD#153	    0.2068	$metal3_conn
Ri83	VDD#153	VDD#154	    0.2068	$metal3_conn
Ri84	VDD#154	VDD#155	    0.2068	$metal3_conn
Ri85	VDD#155	VDD#156	    0.2068	$metal3_conn
Ri86	VDD#156	VDD#157	    0.2068	$metal3_conn
Ri87	VDD#157	VDD#158	    0.2068	$metal3_conn
Ri88	VDD#158	VDD#159	    0.2068	$metal3_conn
Ri89	VDD#159	VDD#160	    0.2068	$metal3_conn
Ri90	VDD#160	VDD#161	    0.2068	$metal3_conn
Ri91	VDD#161	VDD#162	    0.2068	$metal3_conn
Ri92	VDD#162	VDD#163	    0.2068	$metal3_conn
Ri93	VDD#163	VDD#164	    0.2068	$metal3_conn
Ri94	VDD#164	VDD#165	    0.2068	$metal3_conn
Ri95	VDD#165	VDD#166	    0.2068	$metal3_conn
Ri96	VDD#166	VDD#167	    0.2068	$metal3_conn
Ri97	VDD#167	VDD#168	    0.2068	$metal3_conn
Ri98	VDD#168	VDD#169	    0.2068	$metal3_conn
Ri99	VDD#169	VDD#170	    0.2068	$metal3_conn
Ri100	VDD#170	VDD#171	    0.2068	$metal3_conn
Ri101	VDD#171	VDD#172	    0.2068	$metal3_conn
Ri102	VDD#172	VDD#173	    0.2068	$metal3_conn
Ri103	VDD#173	VDD#174	    0.2068	$metal3_conn
Ri104	VDD#174	VDD#175	    0.2068	$metal3_conn
Ri105	VDD#175	VDD#176	    0.2068	$metal3_conn
Ri106	VDD#176	VDD#177	    0.2068	$metal3_conn
Ri107	VDD#177	VDD#178	    0.2068	$metal3_conn
Ri108	VDD#178	VDD#179	    0.2068	$metal3_conn
Ri109	VDD#179	VDD#180	    0.2068	$metal3_conn
Ri110	VDD#180	VDD#181	    0.2068	$metal3_conn
Ri111	VDD#181	VDD#182	    0.2068	$metal3_conn
Ri112	VDD#182	VDD#183	    0.2068	$metal3_conn
Ri113	VDD#183	VDD#184	    0.2068	$metal3_conn
Ri114	VDD#184	VDD#185	    0.2068	$metal3_conn
Ri115	VDD#185	VDD#186	    0.2068	$metal3_conn
Ri116	VDD#186	VDD#187	    0.2068	$metal3_conn
Ri117	VDD#187	VDD#188	    0.2068	$metal3_conn
Ri118	VDD#188	VDD#189	    0.2068	$metal3_conn
Ri119	VDD#189	VDD#190	    0.2068	$metal3_conn
Ri120	VDD#190	VDD#191	    0.2068	$metal3_conn
Ri121	VDD#191	VDD#192	    0.2068	$metal3_conn
Ri122	VDD#192	VDD#193	    0.2068	$metal3_conn
Ri123	VDD#193	VDD#194	    0.2068	$metal3_conn
Ri124	VDD#194	VDD#195	    0.2068	$metal3_conn
Ri125	VDD#195	VDD#196	    0.2068	$metal3_conn
Ri126	VDD#196	VDD#197	    0.2068	$metal3_conn
Ri127	VDD#197	VDD#198	    0.2068	$metal3_conn
Ri128	VDD#198	VDD#200	    0.1378	$metal3_conn
Ri129	VDD	VDD#138	3.954e-02	$metal3_conn
Ri130	VDD#138	VDD#137	    0.2068	$metal3_conn
Ri131	VDD#137	VDD#136	    0.2068	$metal3_conn
Ri132	VDD#136	VDD#135	    0.2068	$metal3_conn
Ri133	VDD#135	VDD#134	    0.2068	$metal3_conn
Ri134	VDD#134	VDD#199	    0.1307	$metal3_conn
Ri135	BLB	BLB#70	    0.3833	$metal3_conn
Ri136	BLB#70	BLB#71	    0.4228	$metal3_conn
Ri137	BLB#71	BLB#72	    0.4228	$metal3_conn
Ri138	BLB#72	BLB#73	    0.4228	$metal3_conn
Ri139	BLB#73	BLB#74	    0.4228	$metal3_conn
Ri140	BLB#74	BLB#75	    0.4228	$metal3_conn
Ri141	BLB#75	BLB#76	    0.4228	$metal3_conn
Ri142	BLB#76	BLB#77	    0.4228	$metal3_conn
Ri143	BLB#77	BLB#78	    0.4228	$metal3_conn
Ri144	BLB#78	BLB#79	    0.4228	$metal3_conn
Ri145	BLB#79	BLB#80	    0.4228	$metal3_conn
Ri146	BLB#80	BLB#81	    0.4228	$metal3_conn
Ri147	BLB#81	BLB#82	    0.4228	$metal3_conn
Ri148	BLB#82	BLB#83	    0.4228	$metal3_conn
Ri149	BLB#83	BLB#84	    0.4228	$metal3_conn
Ri150	BLB#84	BLB#85	    0.4228	$metal3_conn
Ri151	BLB#85	BLB#86	    0.4228	$metal3_conn
Ri152	BLB#86	BLB#87	    0.4228	$metal3_conn
Ri153	BLB#87	BLB#88	    0.4228	$metal3_conn
Ri154	BLB#88	BLB#89	    0.4228	$metal3_conn
Ri155	BLB#89	BLB#90	    0.4228	$metal3_conn
Ri156	BLB#90	BLB#91	    0.4228	$metal3_conn
Ri157	BLB#91	BLB#92	    0.4228	$metal3_conn
Ri158	BLB#92	BLB#93	    0.4228	$metal3_conn
Ri159	BLB#93	BLB#94	    0.4228	$metal3_conn
Ri160	BLB#94	BLB#95	    0.4228	$metal3_conn
Ri161	BLB#95	BLB#96	    0.4228	$metal3_conn
Ri162	BLB#96	BLB#97	    0.4228	$metal3_conn
Ri163	BLB#97	BLB#98	    0.4228	$metal3_conn
Ri164	BLB#98	BLB#99	    0.4324	$metal3_conn
Ri165	BLB	BLB#69	3.954e-02	$metal3_conn
Ri166	BLB#69	BLB#68	    0.4228	$metal3_conn
Ri167	BLB#68	BLB#67	    0.4253	$metal3_conn
Ri168	VSS#70	VSS#173	    7.0179	$metal3_conn
Ri169	VSS#173	VSS#174	    0.4228	$metal3_conn
Ri170	VSS#174	VSS#175	    0.4228	$metal3_conn
Ri171	VSS#175	VSS#176	    0.4228	$metal3_conn
Ri172	VSS#176	VSS#177	    0.4228	$metal3_conn
Ri173	VSS#177	VSS#178	    0.4228	$metal3_conn
Ri174	VSS#178	VSS#179	    0.4228	$metal3_conn
Ri175	VSS#179	VSS#180	    0.4228	$metal3_conn
Ri176	VSS#180	VSS#181	    0.4228	$metal3_conn
Ri177	VSS#181	VSS#182	    0.4228	$metal3_conn
Ri178	VSS#182	VSS#183	    0.4228	$metal3_conn
Ri179	VSS#183	VSS#184	    0.4228	$metal3_conn
Ri180	VSS#184	VSS#185	    0.4228	$metal3_conn
Ri181	VSS#185	VSS#186	    0.4228	$metal3_conn
Ri182	VSS#186	VSS#187	    0.4228	$metal3_conn
Ri183	VSS#187	VSS#188	    0.4228	$metal3_conn
Ri184	VSS#188	VSS#189	    0.4228	$metal3_conn
Ri185	VSS#189	VSS#190	    0.4228	$metal3_conn
Ri186	VSS#190	VSS#191	    0.4228	$metal3_conn
Ri187	VSS#191	VSS#192	    0.4228	$metal3_conn
Ri188	VSS#192	VSS#193	    0.4228	$metal3_conn
Ri189	VSS#193	VSS#194	    0.4228	$metal3_conn
Ri190	VSS#194	VSS#195	    0.4228	$metal3_conn
Ri191	VSS#195	VSS#196	    0.4228	$metal3_conn
Ri192	VSS#196	VSS#197	    0.4228	$metal3_conn
Ri193	VSS#197	VSS#198	    0.4228	$metal3_conn
Ri194	VSS#198	VSS#199	    0.4228	$metal3_conn
Ri195	VSS#199	VSS#200	    0.4228	$metal3_conn
Ri196	VSS#200	VSS#201	    0.4228	$metal3_conn
Ri197	VSS#201	VSS#202	    0.4228	$metal3_conn
Ri198	VSS#202	VSS#203	    0.4228	$metal3_conn
Ri199	VSS#203	VSS#204	    0.4228	$metal3_conn
Ri200	VSS#204	VSS#71	    7.0179	$metal3_conn
*
*       CAPACITOR CARDS
*
*
C1	VDD	VSS	1.50898e-17	$cmodel
C2	WL<0>	VSS	1.14737e-17	$cmodel
C3	WL<10>	VSS	1.14609e-17	$cmodel
C4	WL<11>	VSS	1.14609e-17	$cmodel
C5	WL<12>	VSS	1.14609e-17	$cmodel
C6	WL<13>	VSS	1.14609e-17	$cmodel
C7	WL<14>	VSS	1.14609e-17	$cmodel
C8	WL<15>	VSS	1.14609e-17	$cmodel
C9	WL<16>	VSS	1.14609e-17	$cmodel
C10	WL<17>	VSS	1.14609e-17	$cmodel
C11	WL<18>	VSS	1.14609e-17	$cmodel
C12	WL<19>	VSS	1.14609e-17	$cmodel
C13	WL<1>	VSS	1.14609e-17	$cmodel
C14	WL<20>	VSS	1.14609e-17	$cmodel
C15	WL<21>	VSS	1.14609e-17	$cmodel
C16	WL<22>	VSS	1.14609e-17	$cmodel
C17	WL<23>	VSS	1.14609e-17	$cmodel
C18	WL<24>	VSS	1.14609e-17	$cmodel
C19	WL<25>	VSS	1.14609e-17	$cmodel
C20	WL<26>	VSS	1.14609e-17	$cmodel
C21	WL<27>	VSS	1.14609e-17	$cmodel
C22	WL<28>	VSS	1.14609e-17	$cmodel
C23	WL<29>	VSS	1.14609e-17	$cmodel
C24	WL<2>	VSS	1.14609e-17	$cmodel
C25	WL<30>	VSS	1.14609e-17	$cmodel
C26	WL<31>	VSS	1.14609e-17	$cmodel
C27	WL<32>	VSS	1.14609e-17	$cmodel
C28	WL<33>	VSS	1.14609e-17	$cmodel
C29	WL<34>	VSS	1.14609e-17	$cmodel
C30	WL<35>	VSS	1.14609e-17	$cmodel
C31	WL<36>	VSS	1.14609e-17	$cmodel
C32	WL<37>	VSS	1.14609e-17	$cmodel
C33	WL<38>	VSS	1.14609e-17	$cmodel
C34	WL<39>	VSS	1.14609e-17	$cmodel
C35	WL<3>	VSS	1.14609e-17	$cmodel
C36	WL<40>	VSS	1.14609e-17	$cmodel
C37	WL<41>	VSS	1.14609e-17	$cmodel
C38	WL<42>	VSS	1.14609e-17	$cmodel
C39	WL<43>	VSS	1.14609e-17	$cmodel
C40	WL<44>	VSS	1.14609e-17	$cmodel
C41	WL<45>	VSS	1.14609e-17	$cmodel
C42	WL<46>	VSS	1.14609e-17	$cmodel
C43	WL<47>	VSS	1.14609e-17	$cmodel
C44	WL<48>	VSS	1.14609e-17	$cmodel
C45	WL<49>	VSS	1.14609e-17	$cmodel
C46	WL<4>	VSS	1.14609e-17	$cmodel
C47	WL<50>	VSS	1.14609e-17	$cmodel
C48	WL<51>	VSS	1.14609e-17	$cmodel
C49	WL<52>	VSS	1.14609e-17	$cmodel
C50	WL<53>	VSS	1.14609e-17	$cmodel
C51	WL<54>	VSS	1.14609e-17	$cmodel
C52	WL<55>	VSS	1.14609e-17	$cmodel
C53	WL<56>	VSS	1.14609e-17	$cmodel
C54	WL<57>	VSS	1.14609e-17	$cmodel
C55	WL<58>	VSS	1.14609e-17	$cmodel
C56	WL<59>	VSS	1.14609e-17	$cmodel
C57	WL<5>	VSS	1.14609e-17	$cmodel
C58	WL<60>	VSS	1.14609e-17	$cmodel
C59	WL<61>	VSS	1.14609e-17	$cmodel
C60	WL<62>	VSS	1.14609e-17	$cmodel
C61	WL<63>	VSS	1.14737e-17	$cmodel
C62	WL<6>	VSS	1.14609e-17	$cmodel
C63	WL<7>	VSS	1.14609e-17	$cmodel
C64	WL<8>	VSS	1.14609e-17	$cmodel
C65	WL<9>	VSS	1.14609e-17	$cmodel
C66	BL	VSS	4.31209e-17	$cmodel
C67	BLB	VSS	4.18181e-17	$cmodel
C68	I0<3>/I0<3>/I0<3>/QB	VSS	7.86664e-17	$cmodel
C69	I0<3>/I0<3>/I0<3>/Q	VSS	5.08449e-17	$cmodel
C70	I0<3>/I0<3>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C71	I0<3>/I0<3>/I0<1>/Q	VSS	5.04218e-17	$cmodel
C72	I0<3>/I0<3>/I0<2>/QB	VSS	2.63669e-17	$cmodel
C73	I0<3>/I0<3>/I0<2>/Q	VSS	4.99187e-17	$cmodel
C74	I0<3>/I0<3>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C75	I0<3>/I0<3>/I0<0>/Q	VSS	5.00247e-17	$cmodel
C76	I0<3>/I0<2>/I0<3>/QB	VSS	8.25233e-17	$cmodel
C77	I0<3>/I0<2>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C78	I0<3>/I0<2>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C79	I0<3>/I0<2>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C80	I0<3>/I0<2>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C81	I0<3>/I0<2>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C82	I0<3>/I0<2>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C83	I0<3>/I0<2>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C84	I0<3>/I0<1>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C85	I0<3>/I0<1>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C86	I0<3>/I0<1>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C87	I0<3>/I0<1>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C88	I0<3>/I0<1>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C89	I0<3>/I0<1>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C90	I0<3>/I0<1>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C91	I0<3>/I0<1>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C92	I0<3>/I0<0>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C93	I0<3>/I0<0>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C94	I0<3>/I0<0>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C95	I0<3>/I0<0>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C96	I0<3>/I0<0>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C97	I0<3>/I0<0>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C98	I0<3>/I0<0>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C99	I0<3>/I0<0>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C100	I0<2>/I0<3>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C101	I0<2>/I0<3>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C102	I0<2>/I0<3>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C103	I0<2>/I0<3>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C104	I0<2>/I0<3>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C105	I0<2>/I0<3>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C106	I0<2>/I0<3>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C107	I0<2>/I0<3>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C108	I0<2>/I0<2>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C109	I0<2>/I0<2>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C110	I0<2>/I0<2>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C111	I0<2>/I0<2>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C112	I0<2>/I0<2>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C113	I0<2>/I0<2>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C114	I0<2>/I0<2>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C115	I0<2>/I0<2>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C116	I0<2>/I0<1>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C117	I0<2>/I0<1>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C118	I0<2>/I0<1>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C119	I0<2>/I0<1>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C120	I0<2>/I0<1>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C121	I0<2>/I0<1>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C122	I0<2>/I0<1>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C123	I0<2>/I0<1>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C124	I0<2>/I0<0>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C125	I0<2>/I0<0>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C126	I0<2>/I0<0>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C127	I0<2>/I0<0>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C128	I0<2>/I0<0>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C129	I0<2>/I0<0>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C130	I0<2>/I0<0>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C131	I0<2>/I0<0>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C132	I0<1>/I0<3>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C133	I0<1>/I0<3>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C134	I0<1>/I0<3>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C135	I0<1>/I0<3>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C136	I0<1>/I0<3>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C137	I0<1>/I0<3>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C138	I0<1>/I0<3>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C139	I0<1>/I0<3>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C140	I0<1>/I0<2>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C141	I0<1>/I0<2>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C142	I0<1>/I0<2>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C143	I0<1>/I0<2>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C144	I0<1>/I0<2>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C145	I0<1>/I0<2>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C146	I0<1>/I0<2>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C147	I0<1>/I0<2>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C148	I0<1>/I0<1>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C149	I0<1>/I0<1>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C150	I0<1>/I0<1>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C151	I0<1>/I0<1>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C152	I0<1>/I0<1>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C153	I0<1>/I0<1>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C154	I0<1>/I0<1>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C155	I0<1>/I0<1>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C156	I0<1>/I0<0>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C157	I0<1>/I0<0>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C158	I0<1>/I0<0>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C159	I0<1>/I0<0>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C160	I0<1>/I0<0>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C161	I0<1>/I0<0>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C162	I0<1>/I0<0>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C163	I0<1>/I0<0>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C164	I0<0>/I0<3>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C165	I0<0>/I0<3>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C166	I0<0>/I0<3>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C167	I0<0>/I0<3>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C168	I0<0>/I0<3>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C169	I0<0>/I0<3>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C170	I0<0>/I0<3>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C171	I0<0>/I0<3>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C172	I0<0>/I0<2>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C173	I0<0>/I0<2>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C174	I0<0>/I0<2>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C175	I0<0>/I0<2>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C176	I0<0>/I0<2>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C177	I0<0>/I0<2>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C178	I0<0>/I0<2>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C179	I0<0>/I0<2>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C180	I0<0>/I0<1>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C181	I0<0>/I0<1>/I0<3>/Q	VSS	5.04274e-17	$cmodel
C182	I0<0>/I0<1>/I0<1>/QB	VSS	8.24687e-17	$cmodel
C183	I0<0>/I0<1>/I0<1>/Q	VSS	5.04274e-17	$cmodel
C184	I0<0>/I0<1>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C185	I0<0>/I0<1>/I0<2>/Q	VSS	5.00361e-17	$cmodel
C186	I0<0>/I0<1>/I0<0>/QB	VSS	2.6367e-17	$cmodel
C187	I0<0>/I0<1>/I0<0>/Q	VSS	5.00361e-17	$cmodel
C188	I0<0>/I0<0>/I0<3>/QB	VSS	8.24687e-17	$cmodel
C189	I0<0>/I0<0>/I0<3>/Q	VSS	5.04159e-17	$cmodel
C190	I0<0>/I0<0>/I0<1>/QB	VSS	8.25184e-17	$cmodel
C191	I0<0>/I0<0>/I0<1>/Q	VSS	5.03099e-17	$cmodel
C192	I0<0>/I0<0>/I0<2>/QB	VSS	2.6367e-17	$cmodel
C193	I0<0>/I0<0>/I0<2>/Q	VSS	5.00306e-17	$cmodel
C194	I0<0>/I0<0>/I0<0>/QB	VSS	1.98832e-17	$cmodel
C195	I0<0>/I0<0>/I0<0>/Q	VSS	5.04793e-17	$cmodel
C196	I0<3>/I0<3>/I0<3>/Q#2	VSS	2.75117e-17	$cmodel
C197	I0<3>/I0<3>/I0<2>/Q#2	VSS	2.66779e-17	$cmodel
C198	I0<3>/I0<3>/I0<1>/Q#2	VSS	2.64885e-17	$cmodel
C199	I0<3>/I0<3>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C200	I0<3>/I0<2>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C201	I0<3>/I0<2>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C202	I0<3>/I0<2>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C203	I0<3>/I0<2>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C204	I0<3>/I0<1>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C205	I0<3>/I0<1>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C206	I0<3>/I0<1>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C207	I0<3>/I0<1>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C208	I0<3>/I0<0>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C209	I0<3>/I0<0>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C210	I0<3>/I0<0>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C211	I0<3>/I0<0>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C212	I0<2>/I0<3>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C213	I0<2>/I0<3>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C214	I0<2>/I0<3>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C215	I0<2>/I0<3>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C216	I0<2>/I0<2>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C217	I0<2>/I0<2>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C218	I0<2>/I0<2>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C219	I0<2>/I0<2>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C220	I0<2>/I0<1>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C221	I0<2>/I0<1>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C222	I0<2>/I0<1>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C223	I0<2>/I0<1>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C224	I0<2>/I0<0>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C225	I0<2>/I0<0>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C226	I0<2>/I0<0>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C227	I0<2>/I0<0>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C228	I0<1>/I0<3>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C229	I0<1>/I0<3>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C230	I0<1>/I0<3>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C231	I0<1>/I0<3>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C232	I0<1>/I0<2>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C233	I0<1>/I0<2>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C234	I0<1>/I0<2>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C235	I0<1>/I0<2>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C236	I0<1>/I0<1>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C237	I0<1>/I0<1>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C238	I0<1>/I0<1>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C239	I0<1>/I0<1>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C240	I0<1>/I0<0>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C241	I0<1>/I0<0>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C242	I0<1>/I0<0>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C243	I0<1>/I0<0>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C244	I0<0>/I0<3>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C245	I0<0>/I0<3>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C246	I0<0>/I0<3>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C247	I0<0>/I0<3>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C248	I0<0>/I0<2>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C249	I0<0>/I0<2>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C250	I0<0>/I0<2>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C251	I0<0>/I0<2>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C252	I0<0>/I0<1>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C253	I0<0>/I0<1>/I0<2>/Q#2	VSS	2.64799e-17	$cmodel
C254	I0<0>/I0<1>/I0<1>/Q#2	VSS	2.64799e-17	$cmodel
C255	I0<0>/I0<1>/I0<0>/Q#2	VSS	2.64799e-17	$cmodel
C256	I0<0>/I0<0>/I0<3>/Q#2	VSS	2.64799e-17	$cmodel
C257	I0<0>/I0<0>/I0<2>/Q#2	VSS	2.64885e-17	$cmodel
C258	I0<0>/I0<0>/I0<1>/Q#2	VSS	2.66779e-17	$cmodel
C259	I0<0>/I0<0>/I0<0>/Q#2	VSS	2.75117e-17	$cmodel
C260	I0<3>/I0<3>/I0<3>/QB#2	VSS	1.99934e-17	$cmodel
C261	I0<3>/I0<3>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C262	I0<3>/I0<2>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C263	I0<3>/I0<2>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C264	I0<3>/I0<1>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C265	I0<3>/I0<1>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C266	I0<3>/I0<0>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C267	I0<3>/I0<0>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C268	I0<2>/I0<3>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C269	I0<2>/I0<3>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C270	I0<2>/I0<2>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C271	I0<2>/I0<2>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C272	I0<2>/I0<1>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C273	I0<2>/I0<1>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C274	I0<2>/I0<0>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C275	I0<2>/I0<0>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C276	I0<1>/I0<3>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C277	I0<1>/I0<3>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C278	I0<1>/I0<2>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C279	I0<1>/I0<2>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C280	I0<1>/I0<1>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C281	I0<1>/I0<1>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C282	I0<1>/I0<0>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C283	I0<1>/I0<0>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C284	I0<0>/I0<3>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C285	I0<0>/I0<3>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C286	I0<0>/I0<2>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C287	I0<0>/I0<2>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C288	I0<0>/I0<1>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C289	I0<0>/I0<1>/I0<1>/QB#2	VSS	2.64668e-17	$cmodel
C290	I0<0>/I0<0>/I0<3>/QB#2	VSS	2.64668e-17	$cmodel
C291	I0<0>/I0<0>/I0<1>/QB#2	VSS	2.64667e-17	$cmodel
C292	WL<63>#3	VSS	2.8946e-17	$cmodel
C293	WL<62>#4	VSS	3.56311e-17	$cmodel
C294	WL<61>#3	VSS	3.5558e-17	$cmodel
C295	WL<60>#4	VSS	3.56311e-17	$cmodel
C296	WL<59>#3	VSS	3.5558e-17	$cmodel
C297	WL<58>#4	VSS	3.56311e-17	$cmodel
C298	WL<57>#3	VSS	3.5558e-17	$cmodel
C299	WL<56>#4	VSS	3.56311e-17	$cmodel
C300	WL<55>#3	VSS	3.5558e-17	$cmodel
C301	WL<54>#4	VSS	3.56311e-17	$cmodel
C302	WL<53>#3	VSS	3.5558e-17	$cmodel
C303	WL<52>#4	VSS	3.56311e-17	$cmodel
C304	WL<51>#3	VSS	3.5558e-17	$cmodel
C305	WL<50>#4	VSS	3.56311e-17	$cmodel
C306	WL<49>#3	VSS	3.5558e-17	$cmodel
C307	WL<48>#4	VSS	3.56311e-17	$cmodel
C308	WL<47>#3	VSS	3.5558e-17	$cmodel
C309	WL<46>#4	VSS	3.56311e-17	$cmodel
C310	WL<45>#3	VSS	3.5558e-17	$cmodel
C311	WL<44>#4	VSS	3.56311e-17	$cmodel
C312	WL<43>#3	VSS	3.5558e-17	$cmodel
C313	WL<42>#4	VSS	3.56311e-17	$cmodel
C314	WL<41>#3	VSS	3.5558e-17	$cmodel
C315	WL<40>#4	VSS	3.56311e-17	$cmodel
C316	WL<39>#3	VSS	3.5558e-17	$cmodel
C317	WL<38>#4	VSS	3.56311e-17	$cmodel
C318	WL<37>#3	VSS	3.5558e-17	$cmodel
C319	WL<36>#4	VSS	3.56311e-17	$cmodel
C320	WL<35>#3	VSS	3.5558e-17	$cmodel
C321	WL<34>#4	VSS	3.56311e-17	$cmodel
C322	WL<33>#3	VSS	3.5558e-17	$cmodel
C323	WL<32>#4	VSS	3.56311e-17	$cmodel
C324	WL<31>#3	VSS	3.5558e-17	$cmodel
C325	WL<30>#4	VSS	3.56311e-17	$cmodel
C326	WL<29>#3	VSS	3.5558e-17	$cmodel
C327	WL<28>#4	VSS	3.56311e-17	$cmodel
C328	WL<27>#3	VSS	3.5558e-17	$cmodel
C329	WL<26>#4	VSS	3.56311e-17	$cmodel
C330	WL<25>#3	VSS	3.5558e-17	$cmodel
C331	WL<24>#4	VSS	3.56311e-17	$cmodel
C332	WL<23>#3	VSS	3.5558e-17	$cmodel
C333	WL<22>#4	VSS	3.56311e-17	$cmodel
C334	WL<21>#3	VSS	3.5558e-17	$cmodel
C335	WL<20>#4	VSS	3.56311e-17	$cmodel
C336	WL<19>#3	VSS	3.5558e-17	$cmodel
C337	WL<18>#4	VSS	3.56311e-17	$cmodel
C338	WL<17>#3	VSS	3.5558e-17	$cmodel
C339	WL<16>#4	VSS	3.56311e-17	$cmodel
C340	WL<15>#3	VSS	3.5558e-17	$cmodel
C341	WL<14>#4	VSS	3.56311e-17	$cmodel
C342	WL<13>#3	VSS	3.5558e-17	$cmodel
C343	WL<12>#4	VSS	3.56311e-17	$cmodel
C344	WL<11>#3	VSS	3.5558e-17	$cmodel
C345	WL<10>#4	VSS	3.56311e-17	$cmodel
C346	WL<9>#3	VSS	3.5558e-17	$cmodel
C347	WL<8>#4	VSS	3.56311e-17	$cmodel
C348	WL<7>#3	VSS	3.5558e-17	$cmodel
C349	WL<6>#4	VSS	3.56311e-17	$cmodel
C350	WL<5>#3	VSS	3.5558e-17	$cmodel
C351	WL<4>#4	VSS	3.56311e-17	$cmodel
C352	WL<3>#3	VSS	3.5558e-17	$cmodel
C353	WL<2>#4	VSS	3.56311e-17	$cmodel
C354	WL<1>#3	VSS	3.5558e-17	$cmodel
C355	WL<0>#4	VSS	2.90062e-17	$cmodel
C356	I0<3>/I0<3>/I0<3>/QB#3	VSS	4.17637e-17	$cmodel
C357	WL<63>#1	VSS	3.57766e-17	$cmodel
C358	WL<62>#1	VSS	3.57147e-17	$cmodel
C359	I0<3>/I0<3>/I0<2>/QB#2	VSS	5.04646e-17	$cmodel
C360	I0<3>/I0<3>/I0<1>/QB#3	VSS	5.04673e-17	$cmodel
C361	WL<61>#1	VSS	3.57385e-17	$cmodel
C362	WL<60>#1	VSS	3.56382e-17	$cmodel
C363	I0<3>/I0<3>/I0<0>/QB#2	VSS	5.05094e-17	$cmodel
C364	I0<3>/I0<2>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C365	WL<59>#1	VSS	3.57385e-17	$cmodel
C366	WL<58>#1	VSS	3.56382e-17	$cmodel
C367	I0<3>/I0<2>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C368	I0<3>/I0<2>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C369	WL<57>#1	VSS	3.57385e-17	$cmodel
C370	WL<56>#1	VSS	3.56382e-17	$cmodel
C371	I0<3>/I0<2>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C372	I0<3>/I0<1>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C373	WL<55>#1	VSS	3.57385e-17	$cmodel
C374	WL<54>#1	VSS	3.56382e-17	$cmodel
C375	I0<3>/I0<1>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C376	I0<3>/I0<1>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C377	WL<53>#1	VSS	3.57385e-17	$cmodel
C378	WL<52>#1	VSS	3.56382e-17	$cmodel
C379	I0<3>/I0<1>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C380	I0<3>/I0<0>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C381	WL<51>#1	VSS	3.57385e-17	$cmodel
C382	WL<50>#1	VSS	3.56382e-17	$cmodel
C383	I0<3>/I0<0>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C384	I0<3>/I0<0>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C385	WL<49>#1	VSS	3.57385e-17	$cmodel
C386	WL<48>#1	VSS	3.56382e-17	$cmodel
C387	I0<3>/I0<0>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C388	I0<2>/I0<3>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C389	WL<47>#1	VSS	3.57385e-17	$cmodel
C390	WL<46>#1	VSS	3.56382e-17	$cmodel
C391	I0<2>/I0<3>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C392	I0<2>/I0<3>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C393	WL<45>#1	VSS	3.57385e-17	$cmodel
C394	WL<44>#1	VSS	3.56382e-17	$cmodel
C395	I0<2>/I0<3>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C396	I0<2>/I0<2>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C397	WL<43>#1	VSS	3.57385e-17	$cmodel
C398	WL<42>#1	VSS	3.56382e-17	$cmodel
C399	I0<2>/I0<2>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C400	I0<2>/I0<2>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C401	WL<41>#1	VSS	3.57385e-17	$cmodel
C402	WL<40>#1	VSS	3.56382e-17	$cmodel
C403	I0<2>/I0<2>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C404	I0<2>/I0<1>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C405	WL<39>#1	VSS	3.57385e-17	$cmodel
C406	WL<38>#1	VSS	3.56382e-17	$cmodel
C407	I0<2>/I0<1>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C408	I0<2>/I0<1>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C409	WL<37>#1	VSS	3.57385e-17	$cmodel
C410	WL<36>#1	VSS	3.56382e-17	$cmodel
C411	I0<2>/I0<1>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C412	I0<2>/I0<0>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C413	WL<35>#1	VSS	3.57385e-17	$cmodel
C414	WL<34>#1	VSS	3.56382e-17	$cmodel
C415	I0<2>/I0<0>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C416	I0<2>/I0<0>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C417	WL<33>#1	VSS	3.57385e-17	$cmodel
C418	WL<32>#1	VSS	3.56382e-17	$cmodel
C419	I0<2>/I0<0>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C420	I0<1>/I0<3>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C421	WL<31>#1	VSS	3.57385e-17	$cmodel
C422	WL<30>#1	VSS	3.56382e-17	$cmodel
C423	I0<1>/I0<3>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C424	I0<1>/I0<3>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C425	WL<29>#1	VSS	3.57385e-17	$cmodel
C426	WL<28>#1	VSS	3.56382e-17	$cmodel
C427	I0<1>/I0<3>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C428	I0<1>/I0<2>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C429	WL<27>#1	VSS	3.57385e-17	$cmodel
C430	WL<26>#1	VSS	3.56382e-17	$cmodel
C431	I0<1>/I0<2>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C432	I0<1>/I0<2>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C433	WL<25>#1	VSS	3.57385e-17	$cmodel
C434	WL<24>#1	VSS	3.56382e-17	$cmodel
C435	I0<1>/I0<2>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C436	I0<1>/I0<1>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C437	WL<23>#1	VSS	3.57385e-17	$cmodel
C438	WL<22>#1	VSS	3.56382e-17	$cmodel
C439	I0<1>/I0<1>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C440	I0<1>/I0<1>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C441	WL<21>#1	VSS	3.57385e-17	$cmodel
C442	WL<20>#1	VSS	3.56382e-17	$cmodel
C443	I0<1>/I0<1>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C444	I0<1>/I0<0>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C445	WL<19>#1	VSS	3.57385e-17	$cmodel
C446	WL<18>#1	VSS	3.56382e-17	$cmodel
C447	I0<1>/I0<0>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C448	I0<1>/I0<0>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C449	WL<17>#1	VSS	3.57385e-17	$cmodel
C450	WL<16>#1	VSS	3.56382e-17	$cmodel
C451	I0<1>/I0<0>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C452	I0<0>/I0<3>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C453	WL<15>#1	VSS	3.57385e-17	$cmodel
C454	WL<14>#1	VSS	3.56382e-17	$cmodel
C455	I0<0>/I0<3>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C456	I0<0>/I0<3>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C457	WL<13>#1	VSS	3.57385e-17	$cmodel
C458	WL<12>#1	VSS	3.56382e-17	$cmodel
C459	I0<0>/I0<3>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C460	I0<0>/I0<2>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C461	WL<11>#1	VSS	3.57385e-17	$cmodel
C462	WL<10>#1	VSS	3.56382e-17	$cmodel
C463	I0<0>/I0<2>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C464	I0<0>/I0<2>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C465	WL<9>#1	VSS	3.57385e-17	$cmodel
C466	WL<8>#1	VSS	3.56382e-17	$cmodel
C467	I0<0>/I0<2>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C468	I0<0>/I0<1>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C469	WL<7>#1	VSS	3.57385e-17	$cmodel
C470	WL<6>#1	VSS	3.56382e-17	$cmodel
C471	I0<0>/I0<1>/I0<2>/QB#2	VSS	5.04765e-17	$cmodel
C472	I0<0>/I0<1>/I0<1>/QB#3	VSS	5.04788e-17	$cmodel
C473	WL<5>#1	VSS	3.57385e-17	$cmodel
C474	WL<4>#1	VSS	3.56382e-17	$cmodel
C475	I0<0>/I0<1>/I0<0>/QB#2	VSS	5.04765e-17	$cmodel
C476	I0<0>/I0<0>/I0<3>/QB#3	VSS	5.04788e-17	$cmodel
C477	WL<3>#1	VSS	3.57385e-17	$cmodel
C478	WL<2>#1	VSS	3.56382e-17	$cmodel
C479	I0<0>/I0<0>/I0<2>/QB#2	VSS	5.0465e-17	$cmodel
C480	I0<0>/I0<0>/I0<1>/QB#3	VSS	5.04669e-17	$cmodel
C481	WL<1>#1	VSS	3.5815e-17	$cmodel
C482	WL<0>#1	VSS	3.56762e-17	$cmodel
C483	I0<0>/I0<0>/I0<0>/QB#2	VSS	4.17614e-17	$cmodel
C484	WL<63>#4	VSS	2.14944e-17	$cmodel
C485	WL<62>#3	VSS	3.84451e-17	$cmodel
C486	WL<61>#4	VSS	3.85064e-17	$cmodel
C487	WL<60>#3	VSS	3.84673e-17	$cmodel
C488	WL<59>#4	VSS	3.8517e-17	$cmodel
C489	WL<58>#3	VSS	3.84673e-17	$cmodel
C490	WL<57>#4	VSS	3.8517e-17	$cmodel
C491	WL<56>#3	VSS	3.84673e-17	$cmodel
C492	WL<55>#4	VSS	3.8517e-17	$cmodel
C493	WL<54>#3	VSS	3.84673e-17	$cmodel
C494	WL<53>#4	VSS	3.8517e-17	$cmodel
C495	WL<52>#3	VSS	3.84673e-17	$cmodel
C496	WL<51>#4	VSS	3.8517e-17	$cmodel
C497	WL<50>#3	VSS	3.84673e-17	$cmodel
C498	WL<49>#4	VSS	3.8517e-17	$cmodel
C499	WL<48>#3	VSS	3.84673e-17	$cmodel
C500	WL<47>#4	VSS	3.8517e-17	$cmodel
C501	WL<46>#3	VSS	3.84673e-17	$cmodel
C502	WL<45>#4	VSS	3.8517e-17	$cmodel
C503	WL<44>#3	VSS	3.84673e-17	$cmodel
C504	WL<43>#4	VSS	3.8517e-17	$cmodel
C505	WL<42>#3	VSS	3.84673e-17	$cmodel
C506	WL<41>#4	VSS	3.8517e-17	$cmodel
C507	WL<40>#3	VSS	3.84673e-17	$cmodel
C508	WL<39>#4	VSS	3.8517e-17	$cmodel
C509	WL<38>#3	VSS	3.84673e-17	$cmodel
C510	WL<37>#4	VSS	3.8517e-17	$cmodel
C511	WL<36>#3	VSS	3.84673e-17	$cmodel
C512	WL<35>#4	VSS	3.8517e-17	$cmodel
C513	WL<34>#3	VSS	3.84673e-17	$cmodel
C514	WL<33>#4	VSS	3.8517e-17	$cmodel
C515	WL<32>#3	VSS	3.84673e-17	$cmodel
C516	WL<31>#4	VSS	3.8517e-17	$cmodel
C517	WL<30>#3	VSS	3.84673e-17	$cmodel
C518	WL<29>#4	VSS	3.8517e-17	$cmodel
C519	WL<28>#3	VSS	3.84673e-17	$cmodel
C520	WL<27>#4	VSS	3.8517e-17	$cmodel
C521	WL<26>#3	VSS	3.84673e-17	$cmodel
C522	WL<25>#4	VSS	3.8517e-17	$cmodel
C523	WL<24>#3	VSS	3.84673e-17	$cmodel
C524	WL<23>#4	VSS	3.8517e-17	$cmodel
C525	WL<22>#3	VSS	3.84673e-17	$cmodel
C526	WL<21>#4	VSS	3.8517e-17	$cmodel
C527	WL<20>#3	VSS	3.84673e-17	$cmodel
C528	WL<19>#4	VSS	3.8517e-17	$cmodel
C529	WL<18>#3	VSS	3.84673e-17	$cmodel
C530	WL<17>#4	VSS	3.8517e-17	$cmodel
C531	WL<16>#3	VSS	3.84673e-17	$cmodel
C532	WL<15>#4	VSS	3.8517e-17	$cmodel
C533	WL<14>#3	VSS	3.84673e-17	$cmodel
C534	WL<13>#4	VSS	3.8517e-17	$cmodel
C535	WL<12>#3	VSS	3.84673e-17	$cmodel
C536	WL<11>#4	VSS	3.8517e-17	$cmodel
C537	WL<10>#3	VSS	3.84673e-17	$cmodel
C538	WL<9>#4	VSS	3.8517e-17	$cmodel
C539	WL<8>#3	VSS	3.84673e-17	$cmodel
C540	WL<7>#4	VSS	3.8517e-17	$cmodel
C541	WL<6>#3	VSS	3.84673e-17	$cmodel
C542	WL<5>#4	VSS	3.8517e-17	$cmodel
C543	WL<4>#3	VSS	3.84673e-17	$cmodel
C544	WL<3>#4	VSS	3.8517e-17	$cmodel
C545	WL<2>#3	VSS	3.84567e-17	$cmodel
C546	WL<1>#4	VSS	3.84948e-17	$cmodel
C547	WL<0>#3	VSS	2.14343e-17	$cmodel
C548	I0<3>/I0<3>/I0<2>/QB#3	VSS	8.25887e-17	$cmodel
C549	I0<3>/I0<3>/I0<0>/QB#3	VSS	8.25362e-17	$cmodel
C550	I0<3>/I0<2>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C551	I0<3>/I0<2>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C552	I0<3>/I0<1>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C553	I0<3>/I0<1>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C554	I0<3>/I0<0>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C555	I0<3>/I0<0>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C556	I0<2>/I0<3>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C557	I0<2>/I0<3>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C558	I0<2>/I0<2>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C559	I0<2>/I0<2>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C560	I0<2>/I0<1>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C561	I0<2>/I0<1>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C562	I0<2>/I0<0>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C563	I0<2>/I0<0>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C564	I0<1>/I0<3>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C565	I0<1>/I0<3>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C566	I0<1>/I0<2>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C567	I0<1>/I0<2>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C568	I0<1>/I0<1>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C569	I0<1>/I0<1>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C570	I0<1>/I0<0>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C571	I0<1>/I0<0>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C572	I0<0>/I0<3>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C573	I0<0>/I0<3>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C574	I0<0>/I0<2>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C575	I0<0>/I0<2>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C576	I0<0>/I0<1>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C577	I0<0>/I0<1>/I0<0>/QB#3	VSS	8.2539e-17	$cmodel
C578	I0<0>/I0<0>/I0<2>/QB#3	VSS	8.2539e-17	$cmodel
C579	I0<0>/I0<0>/I0<0>/QB#3	VSS	7.87721e-17	$cmodel
C580	I0<3>/I0<3>/I0<3>/Q#3	VSS	8.28604e-17	$cmodel
C581	I0<3>/I0<3>/I0<2>/Q#3	VSS	8.14159e-17	$cmodel
C582	I0<3>/I0<3>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C583	I0<3>/I0<3>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C584	I0<3>/I0<2>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C585	I0<3>/I0<2>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C586	I0<3>/I0<2>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C587	I0<3>/I0<2>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C588	I0<3>/I0<1>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C589	I0<3>/I0<1>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C590	I0<3>/I0<1>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C591	I0<3>/I0<1>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C592	I0<3>/I0<0>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C593	I0<3>/I0<0>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C594	I0<3>/I0<0>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C595	I0<3>/I0<0>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C596	I0<2>/I0<3>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C597	I0<2>/I0<3>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C598	I0<2>/I0<3>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C599	I0<2>/I0<3>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C600	I0<2>/I0<2>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C601	I0<2>/I0<2>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C602	I0<2>/I0<2>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C603	I0<2>/I0<2>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C604	I0<2>/I0<1>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C605	I0<2>/I0<1>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C606	I0<2>/I0<1>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C607	I0<2>/I0<1>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C608	I0<2>/I0<0>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C609	I0<2>/I0<0>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C610	I0<2>/I0<0>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C611	I0<2>/I0<0>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C612	I0<1>/I0<3>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C613	I0<1>/I0<3>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C614	I0<1>/I0<3>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C615	I0<1>/I0<3>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C616	I0<1>/I0<2>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C617	I0<1>/I0<2>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C618	I0<1>/I0<2>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C619	I0<1>/I0<2>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C620	I0<1>/I0<1>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C621	I0<1>/I0<1>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C622	I0<1>/I0<1>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C623	I0<1>/I0<1>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C624	I0<1>/I0<0>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C625	I0<1>/I0<0>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C626	I0<1>/I0<0>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C627	I0<1>/I0<0>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C628	I0<0>/I0<3>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C629	I0<0>/I0<3>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C630	I0<0>/I0<3>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C631	I0<0>/I0<3>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C632	I0<0>/I0<2>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C633	I0<0>/I0<2>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C634	I0<0>/I0<2>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C635	I0<0>/I0<2>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C636	I0<0>/I0<1>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C637	I0<0>/I0<1>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C638	I0<0>/I0<1>/I0<1>/Q#3	VSS	8.22957e-17	$cmodel
C639	I0<0>/I0<1>/I0<0>/Q#3	VSS	8.14092e-17	$cmodel
C640	I0<0>/I0<0>/I0<3>/Q#3	VSS	8.22957e-17	$cmodel
C641	I0<0>/I0<0>/I0<2>/Q#3	VSS	8.14092e-17	$cmodel
C642	I0<0>/I0<0>/I0<1>/Q#3	VSS	8.23025e-17	$cmodel
C643	I0<0>/I0<0>/I0<0>/Q#3	VSS	8.19476e-17	$cmodel
C644	WL<63>#2	VSS	3.68093e-17	$cmodel
C645	WL<62>#2	VSS	3.62846e-17	$cmodel
C646	WL<61>#2	VSS	3.62952e-17	$cmodel
C647	WL<60>#2	VSS	3.62952e-17	$cmodel
C648	WL<59>#2	VSS	3.62952e-17	$cmodel
C649	WL<58>#2	VSS	3.62952e-17	$cmodel
C650	WL<57>#2	VSS	3.62952e-17	$cmodel
C651	WL<56>#2	VSS	3.62952e-17	$cmodel
C652	WL<55>#2	VSS	3.62952e-17	$cmodel
C653	WL<54>#2	VSS	3.62952e-17	$cmodel
C654	WL<53>#2	VSS	3.62952e-17	$cmodel
C655	WL<52>#2	VSS	3.62952e-17	$cmodel
C656	WL<51>#2	VSS	3.62952e-17	$cmodel
C657	WL<50>#2	VSS	3.62952e-17	$cmodel
C658	WL<49>#2	VSS	3.62952e-17	$cmodel
C659	WL<48>#2	VSS	3.62952e-17	$cmodel
C660	WL<47>#2	VSS	3.62952e-17	$cmodel
C661	WL<46>#2	VSS	3.62952e-17	$cmodel
C662	WL<45>#2	VSS	3.62952e-17	$cmodel
C663	WL<44>#2	VSS	3.62952e-17	$cmodel
C664	WL<43>#2	VSS	3.62952e-17	$cmodel
C665	WL<42>#2	VSS	3.62952e-17	$cmodel
C666	WL<41>#2	VSS	3.62952e-17	$cmodel
C667	WL<40>#2	VSS	3.62952e-17	$cmodel
C668	WL<39>#2	VSS	3.62952e-17	$cmodel
C669	WL<38>#2	VSS	3.62952e-17	$cmodel
C670	WL<37>#2	VSS	3.62952e-17	$cmodel
C671	WL<36>#2	VSS	3.62952e-17	$cmodel
C672	WL<35>#2	VSS	3.62952e-17	$cmodel
C673	WL<34>#2	VSS	3.62952e-17	$cmodel
C674	WL<33>#2	VSS	3.62952e-17	$cmodel
C675	WL<32>#2	VSS	3.62952e-17	$cmodel
C676	WL<31>#2	VSS	3.62952e-17	$cmodel
C677	WL<30>#2	VSS	3.62952e-17	$cmodel
C678	WL<29>#2	VSS	3.62952e-17	$cmodel
C679	WL<28>#2	VSS	3.62952e-17	$cmodel
C680	WL<27>#2	VSS	3.62952e-17	$cmodel
C681	WL<26>#2	VSS	3.62952e-17	$cmodel
C682	WL<25>#2	VSS	3.62952e-17	$cmodel
C683	WL<24>#2	VSS	3.62952e-17	$cmodel
C684	WL<23>#2	VSS	3.62952e-17	$cmodel
C685	WL<22>#2	VSS	3.62952e-17	$cmodel
C686	WL<21>#2	VSS	3.62952e-17	$cmodel
C687	WL<20>#2	VSS	3.62952e-17	$cmodel
C688	WL<19>#2	VSS	3.62952e-17	$cmodel
C689	WL<18>#2	VSS	3.62952e-17	$cmodel
C690	WL<17>#2	VSS	3.62952e-17	$cmodel
C691	WL<16>#2	VSS	3.62952e-17	$cmodel
C692	WL<15>#2	VSS	3.62952e-17	$cmodel
C693	WL<14>#2	VSS	3.62952e-17	$cmodel
C694	WL<13>#2	VSS	3.62952e-17	$cmodel
C695	WL<12>#2	VSS	3.62952e-17	$cmodel
C696	WL<11>#2	VSS	3.62952e-17	$cmodel
C697	WL<10>#2	VSS	3.62952e-17	$cmodel
C698	WL<9>#2	VSS	3.62952e-17	$cmodel
C699	WL<8>#2	VSS	3.62952e-17	$cmodel
C700	WL<7>#2	VSS	3.62952e-17	$cmodel
C701	WL<6>#2	VSS	3.62952e-17	$cmodel
C702	WL<5>#2	VSS	3.62952e-17	$cmodel
C703	WL<4>#2	VSS	3.62952e-17	$cmodel
C704	WL<3>#2	VSS	3.62952e-17	$cmodel
C705	WL<2>#2	VSS	3.62952e-17	$cmodel
C706	WL<1>#2	VSS	3.62846e-17	$cmodel
C707	WL<0>#2	VSS	3.85101e-17	$cmodel
C708	BLB#67	VSS	1.21339e-16	$cmodel
C709	BLB#68	VSS	1.5061e-16	$cmodel
C710	BLB#69	VSS	5.19025e-17	$cmodel
C711	BLB#70	VSS	1.47905e-16	$cmodel
C712	BLB#71	VSS	1.5061e-16	$cmodel
C713	BLB#72	VSS	9.12921e-17	$cmodel
C714	BLB#73	VSS	1.5061e-16	$cmodel
C715	BLB#74	VSS	1.5061e-16	$cmodel
C716	BLB#75	VSS	1.5061e-16	$cmodel
C717	BLB#76	VSS	9.12921e-17	$cmodel
C718	BLB#77	VSS	1.5061e-16	$cmodel
C719	BLB#78	VSS	9.12921e-17	$cmodel
C720	BLB#79	VSS	1.5061e-16	$cmodel
C721	BLB#80	VSS	9.12921e-17	$cmodel
C722	BLB#81	VSS	1.5061e-16	$cmodel
C723	BLB#82	VSS	1.5061e-16	$cmodel
C724	BLB#83	VSS	1.5061e-16	$cmodel
C725	BLB#84	VSS	9.12921e-17	$cmodel
C726	BLB#85	VSS	1.5061e-16	$cmodel
C727	BLB#86	VSS	9.12921e-17	$cmodel
C728	BLB#87	VSS	1.5061e-16	$cmodel
C729	BLB#88	VSS	9.12921e-17	$cmodel
C730	BLB#89	VSS	1.5061e-16	$cmodel
C731	BLB#90	VSS	9.12921e-17	$cmodel
C732	BLB#91	VSS	1.5061e-16	$cmodel
C733	BLB#92	VSS	9.12921e-17	$cmodel
C734	BLB#93	VSS	1.5061e-16	$cmodel
C735	BLB#94	VSS	9.12921e-17	$cmodel
C736	BLB#95	VSS	1.5061e-16	$cmodel
C737	BLB#96	VSS	9.12921e-17	$cmodel
C738	BLB#97	VSS	1.5061e-16	$cmodel
C739	BLB#98	VSS	1.5061e-16	$cmodel
C740	BLB#99	VSS	1.20875e-16	$cmodel
C741	VDD#199	VSS	1.55933e-17	$cmodel
C742	VDD#134	VSS	2.51155e-17	$cmodel
C743	VDD#135	VSS	3.28389e-17	$cmodel
C744	VDD#136	VSS	9.43794e-17	$cmodel
C745	VDD#137	VSS	3.28389e-17	$cmodel
C746	VDD#138	VSS	2.10559e-17	$cmodel
C747	VDD#139	VSS	3.05988e-17	$cmodel
C748	VDD#140	VSS	9.43794e-17	$cmodel
C749	VDD#141	VSS	9.30793e-17	$cmodel
C750	VDD#142	VSS	3.41955e-17	$cmodel
C751	VDD#143	VSS	3.28389e-17	$cmodel
C752	VDD#144	VSS	3.41955e-17	$cmodel
C753	VDD#145	VSS	3.28389e-17	$cmodel
C754	VDD#146	VSS	3.41955e-17	$cmodel
C755	VDD#147	VSS	3.28389e-17	$cmodel
C756	VDD#148	VSS	3.41955e-17	$cmodel
C757	VDD#149	VSS	9.30793e-17	$cmodel
C758	VDD#150	VSS	9.43794e-17	$cmodel
C759	VDD#151	VSS	3.28389e-17	$cmodel
C760	VDD#152	VSS	9.43794e-17	$cmodel
C761	VDD#153	VSS	3.28389e-17	$cmodel
C762	VDD#154	VSS	9.43794e-17	$cmodel
C763	VDD#155	VSS	3.28389e-17	$cmodel
C764	VDD#156	VSS	9.43794e-17	$cmodel
C765	VDD#157	VSS	3.28389e-17	$cmodel
C766	VDD#158	VSS	9.43794e-17	$cmodel
C767	VDD#159	VSS	3.28389e-17	$cmodel
C768	VDD#160	VSS	9.43794e-17	$cmodel
C769	VDD#161	VSS	3.28389e-17	$cmodel
C770	VDD#162	VSS	9.43794e-17	$cmodel
C771	VDD#163	VSS	3.28389e-17	$cmodel
C772	VDD#164	VSS	9.43794e-17	$cmodel
C773	VDD#165	VSS	9.30793e-17	$cmodel
C774	VDD#166	VSS	9.43794e-17	$cmodel
C775	VDD#167	VSS	3.28389e-17	$cmodel
C776	VDD#168	VSS	9.43794e-17	$cmodel
C777	VDD#169	VSS	3.28389e-17	$cmodel
C778	VDD#170	VSS	9.43794e-17	$cmodel
C779	VDD#171	VSS	3.28389e-17	$cmodel
C780	VDD#172	VSS	9.43794e-17	$cmodel
C781	VDD#173	VSS	3.28389e-17	$cmodel
C782	VDD#174	VSS	9.43794e-17	$cmodel
C783	VDD#175	VSS	3.28389e-17	$cmodel
C784	VDD#176	VSS	9.43794e-17	$cmodel
C785	VDD#177	VSS	3.28389e-17	$cmodel
C786	VDD#178	VSS	9.43794e-17	$cmodel
C787	VDD#179	VSS	3.28389e-17	$cmodel
C788	VDD#180	VSS	9.43794e-17	$cmodel
C789	VDD#181	VSS	3.28389e-17	$cmodel
C790	VDD#182	VSS	9.43794e-17	$cmodel
C791	VDD#183	VSS	3.28389e-17	$cmodel
C792	VDD#184	VSS	9.43794e-17	$cmodel
C793	VDD#185	VSS	3.28389e-17	$cmodel
C794	VDD#186	VSS	9.43794e-17	$cmodel
C795	VDD#187	VSS	3.28389e-17	$cmodel
C796	VDD#188	VSS	9.43794e-17	$cmodel
C797	VDD#189	VSS	3.28389e-17	$cmodel
C798	VDD#190	VSS	9.43794e-17	$cmodel
C799	VDD#191	VSS	3.28389e-17	$cmodel
C800	VDD#192	VSS	9.43794e-17	$cmodel
C801	VDD#193	VSS	3.28389e-17	$cmodel
C802	VDD#194	VSS	9.43794e-17	$cmodel
C803	VDD#195	VSS	3.28389e-17	$cmodel
C804	VDD#196	VSS	9.43794e-17	$cmodel
C805	VDD#197	VSS	9.31763e-17	$cmodel
C806	VDD#198	VSS	5.92693e-17	$cmodel
C807	VDD#200	VSS	1.55933e-17	$cmodel
C808	BL#65	VSS	1.78136e-16	$cmodel
C809	BL#66	VSS	1.36196e-16	$cmodel
C810	BL#67	VSS	6.50138e-17	$cmodel
C811	BL#68	VSS	1.52969e-16	$cmodel
C812	BL#69	VSS	1.52969e-16	$cmodel
C813	BL#70	VSS	9.17148e-17	$cmodel
C814	BL#71	VSS	1.52969e-16	$cmodel
C815	BL#72	VSS	1.52969e-16	$cmodel
C816	BL#73	VSS	1.52969e-16	$cmodel
C817	BL#74	VSS	9.17148e-17	$cmodel
C818	BL#75	VSS	1.52969e-16	$cmodel
C819	BL#76	VSS	9.17148e-17	$cmodel
C820	BL#77	VSS	1.52969e-16	$cmodel
C821	BL#78	VSS	9.17148e-17	$cmodel
C822	BL#79	VSS	1.52969e-16	$cmodel
C823	BL#80	VSS	1.52969e-16	$cmodel
C824	BL#81	VSS	1.52969e-16	$cmodel
C825	BL#82	VSS	9.17148e-17	$cmodel
C826	BL#83	VSS	1.52969e-16	$cmodel
C827	BL#84	VSS	9.17148e-17	$cmodel
C828	BL#85	VSS	1.52969e-16	$cmodel
C829	BL#86	VSS	9.17148e-17	$cmodel
C830	BL#87	VSS	1.52969e-16	$cmodel
C831	BL#88	VSS	9.17148e-17	$cmodel
C832	BL#89	VSS	1.52969e-16	$cmodel
C833	BL#90	VSS	9.17148e-17	$cmodel
C834	BL#91	VSS	1.52969e-16	$cmodel
C835	BL#92	VSS	9.17148e-17	$cmodel
C836	BL#93	VSS	1.52969e-16	$cmodel
C837	BL#94	VSS	9.17148e-17	$cmodel
C838	BL#95	VSS	1.52969e-16	$cmodel
C839	BL#96	VSS	1.78136e-16	$cmodel
C840	WL<63>#6	VSS	1.88603e-16	$cmodel
C841	WL<62>#6	VSS	2.05738e-16	$cmodel
C842	WL<61>#6	VSS	2.05612e-16	$cmodel
C843	WL<60>#6	VSS	2.05665e-16	$cmodel
C844	WL<59>#6	VSS	2.05569e-16	$cmodel
C845	WL<58>#6	VSS	2.05665e-16	$cmodel
C846	WL<57>#6	VSS	2.05674e-16	$cmodel
C847	WL<56>#6	VSS	2.05665e-16	$cmodel
C848	WL<55>#6	VSS	2.05674e-16	$cmodel
C849	WL<54>#6	VSS	2.05665e-16	$cmodel
C850	WL<53>#6	VSS	2.05674e-16	$cmodel
C851	WL<52>#6	VSS	2.05665e-16	$cmodel
C852	WL<51>#6	VSS	2.05674e-16	$cmodel
C853	WL<50>#6	VSS	2.05665e-16	$cmodel
C854	WL<49>#6	VSS	2.05674e-16	$cmodel
C855	WL<48>#6	VSS	2.05665e-16	$cmodel
C856	WL<47>#6	VSS	2.05674e-16	$cmodel
C857	WL<46>#6	VSS	2.05665e-16	$cmodel
C858	WL<45>#6	VSS	2.05674e-16	$cmodel
C859	WL<44>#6	VSS	2.05665e-16	$cmodel
C860	WL<43>#6	VSS	2.05674e-16	$cmodel
C861	WL<42>#6	VSS	2.05665e-16	$cmodel
C862	WL<41>#6	VSS	2.05674e-16	$cmodel
C863	WL<40>#6	VSS	2.05665e-16	$cmodel
C864	WL<39>#6	VSS	2.05674e-16	$cmodel
C865	WL<38>#6	VSS	2.05665e-16	$cmodel
C866	WL<37>#6	VSS	2.05674e-16	$cmodel
C867	WL<36>#6	VSS	2.05665e-16	$cmodel
C868	WL<35>#6	VSS	2.05674e-16	$cmodel
C869	WL<34>#6	VSS	2.05665e-16	$cmodel
C870	WL<33>#6	VSS	2.05674e-16	$cmodel
C871	WL<32>#6	VSS	2.05665e-16	$cmodel
C872	WL<31>#6	VSS	2.05674e-16	$cmodel
C873	WL<30>#6	VSS	2.05665e-16	$cmodel
C874	WL<29>#6	VSS	2.05674e-16	$cmodel
C875	WL<28>#6	VSS	2.05665e-16	$cmodel
C876	WL<27>#6	VSS	2.05674e-16	$cmodel
C877	WL<26>#6	VSS	2.05665e-16	$cmodel
C878	WL<25>#6	VSS	2.05674e-16	$cmodel
C879	WL<24>#6	VSS	2.05665e-16	$cmodel
C880	WL<23>#6	VSS	2.05674e-16	$cmodel
C881	WL<22>#6	VSS	2.05665e-16	$cmodel
C882	WL<21>#6	VSS	2.05674e-16	$cmodel
C883	WL<20>#6	VSS	2.05665e-16	$cmodel
C884	WL<19>#6	VSS	2.05674e-16	$cmodel
C885	WL<18>#6	VSS	2.05665e-16	$cmodel
C886	WL<17>#6	VSS	2.05674e-16	$cmodel
C887	WL<16>#6	VSS	2.05665e-16	$cmodel
C888	WL<15>#6	VSS	2.05674e-16	$cmodel
C889	WL<14>#6	VSS	2.05665e-16	$cmodel
C890	WL<13>#6	VSS	2.05674e-16	$cmodel
C891	WL<12>#6	VSS	2.05665e-16	$cmodel
C892	WL<11>#6	VSS	2.05674e-16	$cmodel
C893	WL<10>#6	VSS	2.05665e-16	$cmodel
C894	WL<9>#6	VSS	2.05674e-16	$cmodel
C895	WL<8>#6	VSS	2.05665e-16	$cmodel
C896	WL<7>#6	VSS	2.05674e-16	$cmodel
C897	WL<6>#6	VSS	2.05665e-16	$cmodel
C898	WL<5>#6	VSS	2.05674e-16	$cmodel
C899	WL<4>#6	VSS	2.05665e-16	$cmodel
C900	WL<3>#6	VSS	2.05674e-16	$cmodel
C901	WL<2>#6	VSS	2.05602e-16	$cmodel
C902	WL<1>#6	VSS	2.05748e-16	$cmodel
C903	WL<0>#6	VSS	1.88765e-16	$cmodel
C904	BLB#2	VSS	4.43073e-17	$cmodel
C905	BLB#4	VSS	5.99813e-17	$cmodel
C906	BLB#6	VSS	1.19299e-16	$cmodel
C907	BLB#8	VSS	5.99813e-17	$cmodel
C908	BLB#10	VSS	5.99813e-17	$cmodel
C909	BLB#12	VSS	1.19299e-16	$cmodel
C910	BLB#14	VSS	5.99813e-17	$cmodel
C911	BLB#16	VSS	5.99813e-17	$cmodel
C912	BLB#18	VSS	5.99813e-17	$cmodel
C913	BLB#20	VSS	1.19299e-16	$cmodel
C914	BLB#22	VSS	5.99813e-17	$cmodel
C915	BLB#24	VSS	1.19299e-16	$cmodel
C916	BLB#26	VSS	5.99813e-17	$cmodel
C917	BLB#28	VSS	1.19299e-16	$cmodel
C918	BLB#30	VSS	5.99813e-17	$cmodel
C919	BLB#32	VSS	5.99813e-17	$cmodel
C920	BLB#34	VSS	5.99813e-17	$cmodel
C921	BLB#36	VSS	1.19299e-16	$cmodel
C922	BLB#38	VSS	5.99813e-17	$cmodel
C923	BLB#40	VSS	1.19299e-16	$cmodel
C924	BLB#42	VSS	5.99813e-17	$cmodel
C925	BLB#44	VSS	1.19299e-16	$cmodel
C926	BLB#46	VSS	5.99813e-17	$cmodel
C927	BLB#48	VSS	1.19299e-16	$cmodel
C928	BLB#50	VSS	5.99813e-17	$cmodel
C929	BLB#52	VSS	1.19299e-16	$cmodel
C930	BLB#54	VSS	5.99813e-17	$cmodel
C931	BLB#56	VSS	1.19299e-16	$cmodel
C932	BLB#58	VSS	5.99813e-17	$cmodel
C933	BLB#60	VSS	1.19299e-16	$cmodel
C934	BLB#62	VSS	5.99813e-17	$cmodel
C935	BLB#64	VSS	5.99813e-17	$cmodel
C936	BLB#66	VSS	4.43073e-17	$cmodel
C937	VDD#67	VSS	3.47012e-16	$cmodel
C938	VDD#1	VSS	6.67564e-17	$cmodel
C939	VDD#71	VSS	1.21664e-16	$cmodel
C940	VDD#3	VSS	6.08023e-17	$cmodel
C941	VDD#73	VSS	1.21342e-16	$cmodel
C942	VDD#5	VSS	1.20987e-16	$cmodel
C943	VDD#75	VSS	1.21342e-16	$cmodel
C944	VDD#7	VSS	6.08023e-17	$cmodel
C945	VDD#77	VSS	6.11017e-17	$cmodel
C946	VDD#9	VSS	1.20986e-16	$cmodel
C947	VDD#79	VSS	1.21342e-16	$cmodel
C948	VDD#11	VSS	1.20986e-16	$cmodel
C949	VDD#81	VSS	1.21342e-16	$cmodel
C950	VDD#13	VSS	1.20986e-16	$cmodel
C951	VDD#83	VSS	1.21342e-16	$cmodel
C952	VDD#15	VSS	1.20986e-16	$cmodel
C953	VDD#85	VSS	6.11017e-17	$cmodel
C954	VDD#17	VSS	6.08023e-17	$cmodel
C955	VDD#87	VSS	1.21342e-16	$cmodel
C956	VDD#19	VSS	6.08023e-17	$cmodel
C957	VDD#89	VSS	1.21342e-16	$cmodel
C958	VDD#21	VSS	6.08023e-17	$cmodel
C959	VDD#91	VSS	1.21342e-16	$cmodel
C960	VDD#23	VSS	6.08023e-17	$cmodel
C961	VDD#93	VSS	1.21342e-16	$cmodel
C962	VDD#25	VSS	6.08023e-17	$cmodel
C963	VDD#95	VSS	1.21342e-16	$cmodel
C964	VDD#27	VSS	6.08023e-17	$cmodel
C965	VDD#97	VSS	1.21342e-16	$cmodel
C966	VDD#29	VSS	6.08023e-17	$cmodel
C967	VDD#99	VSS	1.21342e-16	$cmodel
C968	VDD#31	VSS	6.08023e-17	$cmodel
C969	VDD#101	VSS	6.11017e-17	$cmodel
C970	VDD#33	VSS	6.08023e-17	$cmodel
C971	VDD#103	VSS	1.21342e-16	$cmodel
C972	VDD#35	VSS	6.08023e-17	$cmodel
C973	VDD#105	VSS	1.21342e-16	$cmodel
C974	VDD#37	VSS	6.08023e-17	$cmodel
C975	VDD#107	VSS	1.21342e-16	$cmodel
C976	VDD#39	VSS	6.08023e-17	$cmodel
C977	VDD#109	VSS	1.21342e-16	$cmodel
C978	VDD#41	VSS	6.08023e-17	$cmodel
C979	VDD#111	VSS	1.21342e-16	$cmodel
C980	VDD#43	VSS	6.08023e-17	$cmodel
C981	VDD#113	VSS	1.21342e-16	$cmodel
C982	VDD#45	VSS	6.08023e-17	$cmodel
C983	VDD#115	VSS	1.21342e-16	$cmodel
C984	VDD#47	VSS	6.08023e-17	$cmodel
C985	VDD#117	VSS	1.21342e-16	$cmodel
C986	VDD#49	VSS	6.08023e-17	$cmodel
C987	VDD#119	VSS	1.21342e-16	$cmodel
C988	VDD#51	VSS	6.08023e-17	$cmodel
C989	VDD#121	VSS	1.21342e-16	$cmodel
C990	VDD#53	VSS	6.08023e-17	$cmodel
C991	VDD#123	VSS	1.21342e-16	$cmodel
C992	VDD#55	VSS	6.08023e-17	$cmodel
C993	VDD#125	VSS	1.21342e-16	$cmodel
C994	VDD#57	VSS	6.08023e-17	$cmodel
C995	VDD#127	VSS	1.21342e-16	$cmodel
C996	VDD#59	VSS	6.08023e-17	$cmodel
C997	VDD#129	VSS	1.21342e-16	$cmodel
C998	VDD#61	VSS	6.08023e-17	$cmodel
C999	VDD#131	VSS	1.21342e-16	$cmodel
C1000	VDD#63	VSS	6.08023e-17	$cmodel
C1001	VDD#133	VSS	6.13267e-17	$cmodel
C1002	VDD#65	VSS	3.25968e-17	$cmodel
C1003	VDD#69	VSS	3.46777e-16	$cmodel
C1004	BL#2	VSS	6.69504e-17	$cmodel
C1005	BL#4	VSS	6.65929e-17	$cmodel
C1006	BL#6	VSS	1.27847e-16	$cmodel
C1007	BL#8	VSS	6.65929e-17	$cmodel
C1008	BL#10	VSS	6.65929e-17	$cmodel
C1009	BL#12	VSS	1.27847e-16	$cmodel
C1010	BL#14	VSS	6.65929e-17	$cmodel
C1011	BL#16	VSS	6.65929e-17	$cmodel
C1012	BL#18	VSS	6.65929e-17	$cmodel
C1013	BL#20	VSS	1.27847e-16	$cmodel
C1014	BL#22	VSS	6.65929e-17	$cmodel
C1015	BL#24	VSS	1.27847e-16	$cmodel
C1016	BL#26	VSS	6.65929e-17	$cmodel
C1017	BL#28	VSS	1.27847e-16	$cmodel
C1018	BL#30	VSS	6.65929e-17	$cmodel
C1019	BL#32	VSS	6.65929e-17	$cmodel
C1020	BL#34	VSS	6.65929e-17	$cmodel
C1021	BL#36	VSS	1.27847e-16	$cmodel
C1022	BL#38	VSS	6.65929e-17	$cmodel
C1023	BL#40	VSS	1.27847e-16	$cmodel
C1024	BL#42	VSS	6.65929e-17	$cmodel
C1025	BL#44	VSS	1.27847e-16	$cmodel
C1026	BL#46	VSS	6.65929e-17	$cmodel
C1027	BL#48	VSS	1.27847e-16	$cmodel
C1028	BL#50	VSS	6.65929e-17	$cmodel
C1029	BL#52	VSS	1.27847e-16	$cmodel
C1030	BL#54	VSS	6.65929e-17	$cmodel
C1031	BL#56	VSS	1.27847e-16	$cmodel
C1032	BL#58	VSS	6.65929e-17	$cmodel
C1033	BL#60	VSS	1.27847e-16	$cmodel
C1034	BL#62	VSS	6.65929e-17	$cmodel
C1035	BL#64	VSS	6.69504e-17	$cmodel
C1036	WL<63>#5	VSS	6.66564e-17	$cmodel
C1037	WL<62>#5	VSS	6.67349e-17	$cmodel
C1038	WL<61>#5	VSS	6.6517e-17	$cmodel
C1039	WL<60>#5	VSS	6.6517e-17	$cmodel
C1040	WL<59>#5	VSS	6.65411e-17	$cmodel
C1041	WL<58>#5	VSS	6.6517e-17	$cmodel
C1042	WL<57>#5	VSS	6.6517e-17	$cmodel
C1043	WL<56>#5	VSS	6.6517e-17	$cmodel
C1044	WL<55>#5	VSS	6.6517e-17	$cmodel
C1045	WL<54>#5	VSS	6.6517e-17	$cmodel
C1046	WL<53>#5	VSS	6.6517e-17	$cmodel
C1047	WL<52>#5	VSS	6.6517e-17	$cmodel
C1048	WL<51>#5	VSS	6.6517e-17	$cmodel
C1049	WL<50>#5	VSS	6.6517e-17	$cmodel
C1050	WL<49>#5	VSS	6.6517e-17	$cmodel
C1051	WL<48>#5	VSS	6.6517e-17	$cmodel
C1052	WL<47>#5	VSS	6.6517e-17	$cmodel
C1053	WL<46>#5	VSS	6.6517e-17	$cmodel
C1054	WL<45>#5	VSS	6.6517e-17	$cmodel
C1055	WL<44>#5	VSS	6.6517e-17	$cmodel
C1056	WL<43>#5	VSS	6.6517e-17	$cmodel
C1057	WL<42>#5	VSS	6.6517e-17	$cmodel
C1058	WL<41>#5	VSS	6.6517e-17	$cmodel
C1059	WL<40>#5	VSS	6.6517e-17	$cmodel
C1060	WL<39>#5	VSS	6.6517e-17	$cmodel
C1061	WL<38>#5	VSS	6.6517e-17	$cmodel
C1062	WL<37>#5	VSS	6.6517e-17	$cmodel
C1063	WL<36>#5	VSS	6.6517e-17	$cmodel
C1064	WL<35>#5	VSS	6.6517e-17	$cmodel
C1065	WL<34>#5	VSS	6.6517e-17	$cmodel
C1066	WL<33>#5	VSS	6.6517e-17	$cmodel
C1067	WL<32>#5	VSS	6.6517e-17	$cmodel
C1068	WL<31>#5	VSS	6.6517e-17	$cmodel
C1069	WL<30>#5	VSS	6.6517e-17	$cmodel
C1070	WL<29>#5	VSS	6.6517e-17	$cmodel
C1071	WL<28>#5	VSS	6.6517e-17	$cmodel
C1072	WL<27>#5	VSS	6.6517e-17	$cmodel
C1073	WL<26>#5	VSS	6.6517e-17	$cmodel
C1074	WL<25>#5	VSS	6.6517e-17	$cmodel
C1075	WL<24>#5	VSS	6.6517e-17	$cmodel
C1076	WL<23>#5	VSS	6.6517e-17	$cmodel
C1077	WL<22>#5	VSS	6.6517e-17	$cmodel
C1078	WL<21>#5	VSS	6.6517e-17	$cmodel
C1079	WL<20>#5	VSS	6.6517e-17	$cmodel
C1080	WL<19>#5	VSS	6.6517e-17	$cmodel
C1081	WL<18>#5	VSS	6.6517e-17	$cmodel
C1082	WL<17>#5	VSS	6.6517e-17	$cmodel
C1083	WL<16>#5	VSS	6.6517e-17	$cmodel
C1084	WL<15>#5	VSS	6.6517e-17	$cmodel
C1085	WL<14>#5	VSS	6.6517e-17	$cmodel
C1086	WL<13>#5	VSS	6.6517e-17	$cmodel
C1087	WL<12>#5	VSS	6.6517e-17	$cmodel
C1088	WL<11>#5	VSS	6.6517e-17	$cmodel
C1089	WL<10>#5	VSS	6.6517e-17	$cmodel
C1090	WL<9>#5	VSS	6.6517e-17	$cmodel
C1091	WL<8>#5	VSS	6.6517e-17	$cmodel
C1092	WL<7>#5	VSS	6.6517e-17	$cmodel
C1093	WL<6>#5	VSS	6.6517e-17	$cmodel
C1094	WL<5>#5	VSS	6.6517e-17	$cmodel
C1095	WL<4>#5	VSS	6.6517e-17	$cmodel
C1096	WL<3>#5	VSS	6.6517e-17	$cmodel
C1097	WL<2>#5	VSS	6.6517e-17	$cmodel
C1098	WL<1>#5	VSS	6.67349e-17	$cmodel
C1099	WL<0>#5	VSS	6.66564e-17	$cmodel
C1100	VDD#68	VSS	1.22704e-15	$cmodel
C1101	I0<3>/I0<3>/I0<3>/QB#4	VSS	6.11338e-17	$cmodel
C1102	I0<3>/I0<3>/I0<2>/QB#4	VSS	6.01502e-17	$cmodel
C1103	I0<3>/I0<3>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1104	I0<3>/I0<3>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1105	I0<3>/I0<2>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1106	I0<3>/I0<2>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1107	I0<3>/I0<2>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1108	I0<3>/I0<2>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1109	I0<3>/I0<1>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1110	I0<3>/I0<1>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1111	I0<3>/I0<1>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1112	I0<3>/I0<1>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1113	I0<3>/I0<0>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1114	I0<3>/I0<0>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1115	I0<3>/I0<0>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1116	I0<3>/I0<0>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1117	I0<2>/I0<3>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1118	I0<2>/I0<3>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1119	I0<2>/I0<3>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1120	I0<2>/I0<3>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1121	I0<2>/I0<2>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1122	I0<2>/I0<2>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1123	I0<2>/I0<2>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1124	I0<2>/I0<2>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1125	I0<2>/I0<1>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1126	I0<2>/I0<1>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1127	I0<2>/I0<1>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1128	I0<2>/I0<1>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1129	I0<2>/I0<0>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1130	I0<2>/I0<0>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1131	I0<2>/I0<0>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1132	I0<2>/I0<0>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1133	I0<1>/I0<3>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1134	I0<1>/I0<3>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1135	I0<1>/I0<3>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1136	I0<1>/I0<3>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1137	I0<1>/I0<2>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1138	I0<1>/I0<2>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1139	I0<1>/I0<2>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1140	I0<1>/I0<2>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1141	I0<1>/I0<1>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1142	I0<1>/I0<1>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1143	I0<1>/I0<1>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1144	I0<1>/I0<1>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1145	I0<1>/I0<0>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1146	I0<1>/I0<0>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1147	I0<1>/I0<0>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1148	I0<1>/I0<0>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1149	I0<0>/I0<3>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1150	I0<0>/I0<3>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1151	I0<0>/I0<3>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1152	I0<0>/I0<3>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1153	I0<0>/I0<2>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1154	I0<0>/I0<2>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1155	I0<0>/I0<2>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1156	I0<0>/I0<2>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1157	I0<0>/I0<1>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1158	I0<0>/I0<1>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1159	I0<0>/I0<1>/I0<1>/QB#4	VSS	5.98631e-17	$cmodel
C1160	I0<0>/I0<1>/I0<0>/QB#4	VSS	6.01223e-17	$cmodel
C1161	I0<0>/I0<0>/I0<3>/QB#4	VSS	5.98631e-17	$cmodel
C1162	I0<0>/I0<0>/I0<2>/QB#4	VSS	6.01223e-17	$cmodel
C1163	I0<0>/I0<0>/I0<1>/QB#4	VSS	5.9891e-17	$cmodel
C1164	I0<0>/I0<0>/I0<0>/QB#4	VSS	6.14412e-17	$cmodel
C1165	I0<3>/I0<3>/I0<3>/QB#5	VSS	5.70547e-17	$cmodel
C1166	VDD#70	VSS	4.6168e-17	$cmodel
C1167	I0<3>/I0<3>/I0<2>/QB#5	VSS	6.01887e-17	$cmodel
C1168	I0<3>/I0<3>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1169	VDD#72	VSS	4.61336e-17	$cmodel
C1170	I0<3>/I0<3>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1171	I0<3>/I0<2>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1172	VDD#74	VSS	4.61803e-17	$cmodel
C1173	I0<3>/I0<2>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1174	I0<3>/I0<2>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1175	VDD#76	VSS	4.61336e-17	$cmodel
C1176	I0<3>/I0<2>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1177	I0<3>/I0<1>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1178	VDD#78	VSS	4.61336e-17	$cmodel
C1179	I0<3>/I0<1>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1180	I0<3>/I0<1>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1181	VDD#80	VSS	4.61336e-17	$cmodel
C1182	I0<3>/I0<1>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1183	I0<3>/I0<0>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1184	VDD#82	VSS	4.61336e-17	$cmodel
C1185	I0<3>/I0<0>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1186	I0<3>/I0<0>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1187	VDD#84	VSS	4.61336e-17	$cmodel
C1188	I0<3>/I0<0>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1189	I0<2>/I0<3>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1190	VDD#86	VSS	4.61336e-17	$cmodel
C1191	I0<2>/I0<3>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1192	I0<2>/I0<3>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1193	VDD#88	VSS	4.61336e-17	$cmodel
C1194	I0<2>/I0<3>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1195	I0<2>/I0<2>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1196	VDD#90	VSS	4.61336e-17	$cmodel
C1197	I0<2>/I0<2>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1198	I0<2>/I0<2>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1199	VDD#92	VSS	4.61336e-17	$cmodel
C1200	I0<2>/I0<2>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1201	I0<2>/I0<1>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1202	VDD#94	VSS	4.61336e-17	$cmodel
C1203	I0<2>/I0<1>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1204	I0<2>/I0<1>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1205	VDD#96	VSS	4.61336e-17	$cmodel
C1206	I0<2>/I0<1>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1207	I0<2>/I0<0>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1208	VDD#98	VSS	4.61336e-17	$cmodel
C1209	I0<2>/I0<0>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1210	I0<2>/I0<0>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1211	VDD#100	VSS	4.61336e-17	$cmodel
C1212	I0<2>/I0<0>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1213	I0<1>/I0<3>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1214	VDD#102	VSS	4.61336e-17	$cmodel
C1215	I0<1>/I0<3>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1216	I0<1>/I0<3>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1217	VDD#104	VSS	4.61336e-17	$cmodel
C1218	I0<1>/I0<3>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1219	I0<1>/I0<2>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1220	VDD#106	VSS	4.61336e-17	$cmodel
C1221	I0<1>/I0<2>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1222	I0<1>/I0<2>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1223	VDD#108	VSS	4.61336e-17	$cmodel
C1224	I0<1>/I0<2>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1225	I0<1>/I0<1>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1226	VDD#110	VSS	4.61336e-17	$cmodel
C1227	I0<1>/I0<1>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1228	I0<1>/I0<1>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1229	VDD#112	VSS	4.61336e-17	$cmodel
C1230	I0<1>/I0<1>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1231	I0<1>/I0<0>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1232	VDD#114	VSS	4.61336e-17	$cmodel
C1233	I0<1>/I0<0>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1234	I0<1>/I0<0>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1235	VDD#116	VSS	4.61336e-17	$cmodel
C1236	I0<1>/I0<0>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1237	I0<0>/I0<3>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1238	VDD#118	VSS	4.61336e-17	$cmodel
C1239	I0<0>/I0<3>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1240	I0<0>/I0<3>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1241	VDD#120	VSS	4.61336e-17	$cmodel
C1242	I0<0>/I0<3>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1243	I0<0>/I0<2>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1244	VDD#122	VSS	4.61336e-17	$cmodel
C1245	I0<0>/I0<2>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1246	I0<0>/I0<2>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1247	VDD#124	VSS	4.61336e-17	$cmodel
C1248	I0<0>/I0<2>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1249	I0<0>/I0<1>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1250	VDD#126	VSS	4.61336e-17	$cmodel
C1251	I0<0>/I0<1>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1252	I0<0>/I0<1>/I0<1>/QB#5	VSS	6.00461e-17	$cmodel
C1253	VDD#128	VSS	4.61336e-17	$cmodel
C1254	I0<0>/I0<1>/I0<0>/QB#5	VSS	6.00463e-17	$cmodel
C1255	I0<0>/I0<0>/I0<3>/QB#5	VSS	6.00461e-17	$cmodel
C1256	VDD#130	VSS	4.61336e-17	$cmodel
C1257	I0<0>/I0<0>/I0<2>/QB#5	VSS	6.00463e-17	$cmodel
C1258	I0<0>/I0<0>/I0<1>/QB#5	VSS	6.01885e-17	$cmodel
C1259	VDD#132	VSS	4.6168e-17	$cmodel
C1260	I0<0>/I0<0>/I0<0>/QB#5	VSS	5.72465e-17	$cmodel
C1261	VDD#2	VSS	2.84073e-17	$cmodel
C1262	I0<3>/I0<3>/I0<3>/Q#4	VSS	5.17174e-17	$cmodel
C1263	I0<3>/I0<3>/I0<2>/Q#4	VSS	5.85908e-17	$cmodel
C1264	VDD#4	VSS	4.68023e-17	$cmodel
C1265	I0<3>/I0<3>/I0<1>/Q#4	VSS	5.85476e-17	$cmodel
C1266	I0<3>/I0<3>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1267	VDD#6	VSS	4.67538e-17	$cmodel
C1268	I0<3>/I0<2>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1269	I0<3>/I0<2>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1270	VDD#8	VSS	4.675e-17	$cmodel
C1271	I0<3>/I0<2>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1272	I0<3>/I0<2>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1273	VDD#10	VSS	4.675e-17	$cmodel
C1274	I0<3>/I0<1>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1275	I0<3>/I0<1>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1276	VDD#12	VSS	4.675e-17	$cmodel
C1277	I0<3>/I0<1>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1278	I0<3>/I0<1>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1279	VDD#14	VSS	4.675e-17	$cmodel
C1280	I0<3>/I0<0>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1281	I0<3>/I0<0>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1282	VDD#16	VSS	4.675e-17	$cmodel
C1283	I0<3>/I0<0>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1284	I0<3>/I0<0>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1285	VDD#18	VSS	4.675e-17	$cmodel
C1286	I0<2>/I0<3>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1287	I0<2>/I0<3>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1288	VDD#20	VSS	4.675e-17	$cmodel
C1289	I0<2>/I0<3>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1290	I0<2>/I0<3>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1291	VDD#22	VSS	4.675e-17	$cmodel
C1292	I0<2>/I0<2>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1293	I0<2>/I0<2>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1294	VDD#24	VSS	4.675e-17	$cmodel
C1295	I0<2>/I0<2>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1296	I0<2>/I0<2>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1297	VDD#26	VSS	4.675e-17	$cmodel
C1298	I0<2>/I0<1>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1299	I0<2>/I0<1>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1300	VDD#28	VSS	4.675e-17	$cmodel
C1301	I0<2>/I0<1>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1302	I0<2>/I0<1>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1303	VDD#30	VSS	4.675e-17	$cmodel
C1304	I0<2>/I0<0>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1305	I0<2>/I0<0>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1306	VDD#32	VSS	4.675e-17	$cmodel
C1307	I0<2>/I0<0>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1308	I0<2>/I0<0>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1309	VDD#34	VSS	4.675e-17	$cmodel
C1310	I0<1>/I0<3>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1311	I0<1>/I0<3>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1312	VDD#36	VSS	4.675e-17	$cmodel
C1313	I0<1>/I0<3>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1314	I0<1>/I0<3>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1315	VDD#38	VSS	4.675e-17	$cmodel
C1316	I0<1>/I0<2>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1317	I0<1>/I0<2>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1318	VDD#40	VSS	4.675e-17	$cmodel
C1319	I0<1>/I0<2>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1320	I0<1>/I0<2>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1321	VDD#42	VSS	4.675e-17	$cmodel
C1322	I0<1>/I0<1>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1323	I0<1>/I0<1>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1324	VDD#44	VSS	4.675e-17	$cmodel
C1325	I0<1>/I0<1>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1326	I0<1>/I0<1>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1327	VDD#46	VSS	4.675e-17	$cmodel
C1328	I0<1>/I0<0>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1329	I0<1>/I0<0>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1330	VDD#48	VSS	4.675e-17	$cmodel
C1331	I0<1>/I0<0>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1332	I0<1>/I0<0>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1333	VDD#50	VSS	4.675e-17	$cmodel
C1334	I0<0>/I0<3>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1335	I0<0>/I0<3>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1336	VDD#52	VSS	4.675e-17	$cmodel
C1337	I0<0>/I0<3>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1338	I0<0>/I0<3>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1339	VDD#54	VSS	4.675e-17	$cmodel
C1340	I0<0>/I0<2>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1341	I0<0>/I0<2>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1342	VDD#56	VSS	4.675e-17	$cmodel
C1343	I0<0>/I0<2>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1344	I0<0>/I0<2>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1345	VDD#58	VSS	4.675e-17	$cmodel
C1346	I0<0>/I0<1>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1347	I0<0>/I0<1>/I0<2>/Q#4	VSS	5.84786e-17	$cmodel
C1348	VDD#60	VSS	4.675e-17	$cmodel
C1349	I0<0>/I0<1>/I0<1>/Q#4	VSS	5.84786e-17	$cmodel
C1350	I0<0>/I0<1>/I0<0>/Q#4	VSS	5.84786e-17	$cmodel
C1351	VDD#62	VSS	4.675e-17	$cmodel
C1352	I0<0>/I0<0>/I0<3>/Q#4	VSS	5.84786e-17	$cmodel
C1353	I0<0>/I0<0>/I0<2>/Q#4	VSS	5.85476e-17	$cmodel
C1354	VDD#64	VSS	4.68023e-17	$cmodel
C1355	I0<0>/I0<0>/I0<1>/Q#4	VSS	5.85908e-17	$cmodel
C1356	I0<0>/I0<0>/I0<0>/Q#4	VSS	5.2584e-17	$cmodel
C1357	VDD#66	VSS	2.84097e-17	$cmodel
C1358	I0<3>/I0<3>/I0<3>/Q#6	VSS	6.02111e-17	$cmodel
C1359	I0<3>/I0<3>/I0<2>/Q#6	VSS	6.28358e-17	$cmodel
C1360	I0<3>/I0<3>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1361	I0<3>/I0<3>/I0<0>/Q#6	VSS	6.27526e-17	$cmodel
C1362	I0<3>/I0<2>/I0<3>/Q#6	VSS	6.28425e-17	$cmodel
C1363	I0<3>/I0<2>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1364	I0<3>/I0<2>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1365	I0<3>/I0<2>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1366	I0<3>/I0<1>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1367	I0<3>/I0<1>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1368	I0<3>/I0<1>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1369	I0<3>/I0<1>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1370	I0<3>/I0<0>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1371	I0<3>/I0<0>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1372	I0<3>/I0<0>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1373	I0<3>/I0<0>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1374	I0<2>/I0<3>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1375	I0<2>/I0<3>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1376	I0<2>/I0<3>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1377	I0<2>/I0<3>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1378	I0<2>/I0<2>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1379	I0<2>/I0<2>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1380	I0<2>/I0<2>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1381	I0<2>/I0<2>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1382	I0<2>/I0<1>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1383	I0<2>/I0<1>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1384	I0<2>/I0<1>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1385	I0<2>/I0<1>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1386	I0<2>/I0<0>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1387	I0<2>/I0<0>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1388	I0<2>/I0<0>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1389	I0<2>/I0<0>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1390	I0<1>/I0<3>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1391	I0<1>/I0<3>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1392	I0<1>/I0<3>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1393	I0<1>/I0<3>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1394	I0<1>/I0<2>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1395	I0<1>/I0<2>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1396	I0<1>/I0<2>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1397	I0<1>/I0<2>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1398	I0<1>/I0<1>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1399	I0<1>/I0<1>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1400	I0<1>/I0<1>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1401	I0<1>/I0<1>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1402	I0<1>/I0<0>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1403	I0<1>/I0<0>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1404	I0<1>/I0<0>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1405	I0<1>/I0<0>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1406	I0<0>/I0<3>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1407	I0<0>/I0<3>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1408	I0<0>/I0<3>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1409	I0<0>/I0<3>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1410	I0<0>/I0<2>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1411	I0<0>/I0<2>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1412	I0<0>/I0<2>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1413	I0<0>/I0<2>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1414	I0<0>/I0<1>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1415	I0<0>/I0<1>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1416	I0<0>/I0<1>/I0<1>/Q#6	VSS	6.28084e-17	$cmodel
C1417	I0<0>/I0<1>/I0<0>/Q#6	VSS	6.28084e-17	$cmodel
C1418	I0<0>/I0<0>/I0<3>/Q#6	VSS	6.28084e-17	$cmodel
C1419	I0<0>/I0<0>/I0<2>/Q#6	VSS	6.28084e-17	$cmodel
C1420	I0<0>/I0<0>/I0<1>/Q#6	VSS	6.28358e-17	$cmodel
C1421	I0<0>/I0<0>/I0<0>/Q#6	VSS	6.09442e-17	$cmodel
C1422	WL<63>#7	VSS	1.35933e-16	$cmodel
C1423	WL<62>#7	VSS	1.42746e-16	$cmodel
C1424	WL<61>#7	VSS	1.42552e-16	$cmodel
C1425	WL<60>#7	VSS	1.42542e-16	$cmodel
C1426	WL<59>#7	VSS	1.42419e-16	$cmodel
C1427	WL<58>#7	VSS	1.42542e-16	$cmodel
C1428	WL<57>#7	VSS	1.42544e-16	$cmodel
C1429	WL<56>#7	VSS	1.42542e-16	$cmodel
C1430	WL<55>#7	VSS	1.42544e-16	$cmodel
C1431	WL<54>#7	VSS	1.42542e-16	$cmodel
C1432	WL<53>#7	VSS	1.42544e-16	$cmodel
C1433	WL<52>#7	VSS	1.42542e-16	$cmodel
C1434	WL<51>#7	VSS	1.42544e-16	$cmodel
C1435	WL<50>#7	VSS	1.42542e-16	$cmodel
C1436	WL<49>#7	VSS	1.42544e-16	$cmodel
C1437	WL<48>#7	VSS	1.42542e-16	$cmodel
C1438	WL<47>#7	VSS	1.42544e-16	$cmodel
C1439	WL<46>#7	VSS	1.42542e-16	$cmodel
C1440	WL<45>#7	VSS	1.42544e-16	$cmodel
C1441	WL<44>#7	VSS	1.42542e-16	$cmodel
C1442	WL<43>#7	VSS	1.42544e-16	$cmodel
C1443	WL<42>#7	VSS	1.42542e-16	$cmodel
C1444	WL<41>#7	VSS	1.42544e-16	$cmodel
C1445	WL<40>#7	VSS	1.42542e-16	$cmodel
C1446	WL<39>#7	VSS	1.42544e-16	$cmodel
C1447	WL<38>#7	VSS	1.42542e-16	$cmodel
C1448	WL<37>#7	VSS	1.42544e-16	$cmodel
C1449	WL<36>#7	VSS	1.42542e-16	$cmodel
C1450	WL<35>#7	VSS	1.42544e-16	$cmodel
C1451	WL<34>#7	VSS	1.42542e-16	$cmodel
C1452	WL<33>#7	VSS	1.42544e-16	$cmodel
C1453	WL<32>#7	VSS	1.42542e-16	$cmodel
C1454	WL<31>#7	VSS	1.42544e-16	$cmodel
C1455	WL<30>#7	VSS	1.42542e-16	$cmodel
C1456	WL<29>#7	VSS	1.42544e-16	$cmodel
C1457	WL<28>#7	VSS	1.42542e-16	$cmodel
C1458	WL<27>#7	VSS	1.42544e-16	$cmodel
C1459	WL<26>#7	VSS	1.42542e-16	$cmodel
C1460	WL<25>#7	VSS	1.42544e-16	$cmodel
C1461	WL<24>#7	VSS	1.42542e-16	$cmodel
C1462	WL<23>#7	VSS	1.42544e-16	$cmodel
C1463	WL<22>#7	VSS	1.42542e-16	$cmodel
C1464	WL<21>#7	VSS	1.42544e-16	$cmodel
C1465	WL<20>#7	VSS	1.42542e-16	$cmodel
C1466	WL<19>#7	VSS	1.42544e-16	$cmodel
C1467	WL<18>#7	VSS	1.42542e-16	$cmodel
C1468	WL<17>#7	VSS	1.42544e-16	$cmodel
C1469	WL<16>#7	VSS	1.42542e-16	$cmodel
C1470	WL<15>#7	VSS	1.42544e-16	$cmodel
C1471	WL<14>#7	VSS	1.42542e-16	$cmodel
C1472	WL<13>#7	VSS	1.42544e-16	$cmodel
C1473	WL<12>#7	VSS	1.42542e-16	$cmodel
C1474	WL<11>#7	VSS	1.42544e-16	$cmodel
C1475	WL<10>#7	VSS	1.42542e-16	$cmodel
C1476	WL<9>#7	VSS	1.42544e-16	$cmodel
C1477	WL<8>#7	VSS	1.42542e-16	$cmodel
C1478	WL<7>#7	VSS	1.42544e-16	$cmodel
C1479	WL<6>#7	VSS	1.42542e-16	$cmodel
C1480	WL<5>#7	VSS	1.42544e-16	$cmodel
C1481	WL<4>#7	VSS	1.42542e-16	$cmodel
C1482	WL<3>#7	VSS	1.42544e-16	$cmodel
C1483	WL<2>#7	VSS	1.4255e-16	$cmodel
C1484	WL<1>#7	VSS	1.42747e-16	$cmodel
C1485	WL<0>#7	VSS	1.37485e-16	$cmodel
*
*
.ENDS bit_cell_col_64
*

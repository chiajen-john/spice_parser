*
*
*
*                       LINUX           Thu Nov 23 18:02:06 2023
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus - (64-bit)
*  Version        : 19.1.3-s062
*  Build Date     : Tue Jul 23 02:42:20 PDT 2019
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT bit_cell_row_64 VDD VSS WL BL<0> BL<10> BL<11> BL<12> BL<13> BL<14>
+ BL<15> BL<16> BL<17> BL<18> BL<19> BL<1> BL<20> BL<21> BL<22> BL<23> BL<24>
+ BL<25> BL<26> BL<27> BL<28> BL<29> BL<2> BL<30> BL<31> BL<32> BL<33> BL<34>
+ BL<35> BL<36> BL<37> BL<38> BL<39> BL<3> BL<40> BL<41> BL<42> BL<43> BL<44>
+ BL<45> BL<46> BL<47> BL<48> BL<49> BL<4> BL<50> BL<51> BL<52> BL<53> BL<54>
+ BL<55> BL<56> BL<57> BL<58> BL<59> BL<5> BL<60> BL<61> BL<62> BL<63> BL<6>
+ BL<7> BL<8> BL<9> BLB<0> BLB<10> BLB<11> BLB<12> BLB<13> BLB<14> BLB<15>
+ BLB<16> BLB<17> BLB<18> BLB<19> BLB<1> BLB<20> BLB<21> BLB<22> BLB<23> BLB<24>
+ BLB<25> BLB<26> BLB<27> BLB<28> BLB<29> BLB<2> BLB<30> BLB<31> BLB<32> BLB<33>
+ BLB<34> BLB<35> BLB<36> BLB<37> BLB<38> BLB<39> BLB<3> BLB<40> BLB<41> BLB<42>
+ BLB<43> BLB<44> BLB<45> BLB<46> BLB<47> BLB<48> BLB<49> BLB<4> BLB<50> BLB<51>
+ BLB<52> BLB<53> BLB<54> BLB<55> BLB<56> BLB<57> BLB<58> BLB<59> BLB<5> BLB<60>
+ BLB<61> BLB<62> BLB<63> BLB<6> BLB<7> BLB<8> BLB<9>
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MI0<7>/I1<7>/NM0	I0<7>/I1<7>/Q#4	WL#254	BL<63>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<7>/NM2	I0<7>/I1<7>/Q#4	I0<7>/I1<7>/QB	VSS#383
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<7>/NM1	BLB<63>#1	WL#250	I0<7>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<7>/NM3	I0<7>/I1<7>/QB#6	I0<7>/I1<7>/Q#3	VSS#378
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<6>/NM0	I0<7>/I1<6>/Q#4	WL#248	BL<61>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<6>/NM2	I0<7>/I1<6>/Q#4	I0<7>/I1<6>/QB	VSS#376
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<6>/NM1	BLB<61>#1	WL#242	I0<7>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<6>/NM3	I0<7>/I1<6>/QB#6	I0<7>/I1<6>/Q#3	VSS#371
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<5>/NM0	I0<7>/I1<5>/Q#6	WL#246	BL<62>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<5>/NM2	I0<7>/I1<5>/Q#6	I0<7>/I1<5>/QB#2	VSS#374
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<5>/NM1	BLB<62>#1	WL#252	I0<7>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<5>/NM3	I0<7>/I1<5>/QB#4	I0<7>/I1<5>/Q	VSS#380
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<4>/NM0	I0<7>/I1<4>/Q#4	WL#240	BL<59>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<4>/NM2	I0<7>/I1<4>/Q#4	I0<7>/I1<4>/QB	VSS#366
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<4>/NM1	BLB<59>#1	WL#234	I0<7>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<4>/NM3	I0<7>/I1<4>/QB#6	I0<7>/I1<4>/Q#3	VSS#359
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<3>/NM0	I0<7>/I1<3>/Q#6	WL#238	BL<60>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<3>/NM2	I0<7>/I1<3>/Q#6	I0<7>/I1<3>/QB#2	VSS#365
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<3>/NM1	BLB<60>#3	WL#244	I0<7>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<3>/NM3	I0<7>/I1<3>/QB#4	I0<7>/I1<3>/Q	VSS#372
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<2>/NM0	I0<7>/I1<2>/Q#4	WL#232	BL<57>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<2>/NM2	I0<7>/I1<2>/Q#4	I0<7>/I1<2>/QB	VSS#354
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<2>/NM1	BLB<57>#1	WL#226	I0<7>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<2>/NM3	I0<7>/I1<2>/QB#6	I0<7>/I1<2>/Q#3	VSS#347
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<1>/NM0	I0<7>/I1<1>/Q#6	WL#230	BL<58>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<1>/NM2	I0<7>/I1<1>/Q#6	I0<7>/I1<1>/QB#2	VSS#353
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<1>/NM1	BLB<58>#3	WL#236	I0<7>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<1>/NM3	I0<7>/I1<1>/QB#4	I0<7>/I1<1>/Q	VSS#360
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<0>/NM0	I0<7>/I1<0>/Q#6	WL#222	BL<56>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<0>/NM2	I0<7>/I1<0>/Q#6	I0<7>/I1<0>/QB#2	VSS#341
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<0>/NM1	BLB<56>#3	WL#228	I0<7>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<7>/I1<0>/NM3	I0<7>/I1<0>/QB#4	I0<7>/I1<0>/Q	VSS#348
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<7>/NM0	I0<6>/I1<7>/Q#4	WL#224	BL<55>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<7>/NM2	I0<6>/I1<7>/Q#4	I0<6>/I1<7>/QB	VSS#342
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<7>/NM1	BLB<55>#1	WL#218	I0<6>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<7>/NM3	I0<6>/I1<7>/QB#6	I0<6>/I1<7>/Q#3	VSS#335
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<6>/NM0	I0<6>/I1<6>/Q#4	WL#216	BL<53>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<6>/NM2	I0<6>/I1<6>/Q#4	I0<6>/I1<6>/QB	VSS#330
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<6>/NM1	BLB<53>#1	WL#210	I0<6>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<6>/NM3	I0<6>/I1<6>/QB#6	I0<6>/I1<6>/Q#3	VSS#323
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<5>/NM0	I0<6>/I1<5>/Q#6	WL#214	BL<54>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<5>/NM2	I0<6>/I1<5>/Q#6	I0<6>/I1<5>/QB#2	VSS#329
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<5>/NM1	BLB<54>#3	WL#220	I0<6>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<5>/NM3	I0<6>/I1<5>/QB#4	I0<6>/I1<5>/Q	VSS#336
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<4>/NM0	I0<6>/I1<4>/Q#4	WL#208	BL<51>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<4>/NM2	I0<6>/I1<4>/Q#4	I0<6>/I1<4>/QB	VSS#318
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<4>/NM1	BLB<51>#1	WL#202	I0<6>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<4>/NM3	I0<6>/I1<4>/QB#6	I0<6>/I1<4>/Q#3	VSS#311
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<3>/NM0	I0<6>/I1<3>/Q#6	WL#206	BL<52>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<3>/NM2	I0<6>/I1<3>/Q#6	I0<6>/I1<3>/QB#2	VSS#317
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<3>/NM1	BLB<52>#3	WL#212	I0<6>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<3>/NM3	I0<6>/I1<3>/QB#4	I0<6>/I1<3>/Q	VSS#324
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<2>/NM0	I0<6>/I1<2>/Q#4	WL#200	BL<49>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<2>/NM2	I0<6>/I1<2>/Q#4	I0<6>/I1<2>/QB	VSS#306
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<2>/NM1	BLB<49>#1	WL#194	I0<6>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<2>/NM3	I0<6>/I1<2>/QB#6	I0<6>/I1<2>/Q#3	VSS#299
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<1>/NM0	I0<6>/I1<1>/Q#6	WL#198	BL<50>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<1>/NM2	I0<6>/I1<1>/Q#6	I0<6>/I1<1>/QB#2	VSS#305
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<1>/NM1	BLB<50>#3	WL#204	I0<6>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<1>/NM3	I0<6>/I1<1>/QB#4	I0<6>/I1<1>/Q	VSS#312
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<0>/NM0	I0<6>/I1<0>/Q#6	WL#190	BL<48>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<0>/NM2	I0<6>/I1<0>/Q#6	I0<6>/I1<0>/QB#2	VSS#293
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<6>/I1<0>/NM1	BLB<48>#3	WL#196	I0<6>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<6>/I1<0>/NM3	I0<6>/I1<0>/QB#4	I0<6>/I1<0>/Q	VSS#300
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<7>/NM0	I0<5>/I1<7>/Q#4	WL#192	BL<47>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<7>/NM2	I0<5>/I1<7>/Q#4	I0<5>/I1<7>/QB	VSS#294
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<7>/NM1	BLB<47>#1	WL#186	I0<5>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<7>/NM3	I0<5>/I1<7>/QB#6	I0<5>/I1<7>/Q#3	VSS#287
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<6>/NM0	I0<5>/I1<6>/Q#4	WL#184	BL<45>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<6>/NM2	I0<5>/I1<6>/Q#4	I0<5>/I1<6>/QB	VSS#282
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<6>/NM1	BLB<45>#1	WL#178	I0<5>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<6>/NM3	I0<5>/I1<6>/QB#6	I0<5>/I1<6>/Q#3	VSS#275
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<5>/NM0	I0<5>/I1<5>/Q#6	WL#182	BL<46>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<5>/NM2	I0<5>/I1<5>/Q#6	I0<5>/I1<5>/QB#2	VSS#281
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<5>/NM1	BLB<46>#3	WL#188	I0<5>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<5>/NM3	I0<5>/I1<5>/QB#4	I0<5>/I1<5>/Q	VSS#288
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<4>/NM0	I0<5>/I1<4>/Q#4	WL#176	BL<43>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<4>/NM2	I0<5>/I1<4>/Q#4	I0<5>/I1<4>/QB	VSS#270
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<4>/NM1	BLB<43>#1	WL#170	I0<5>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<4>/NM3	I0<5>/I1<4>/QB#6	I0<5>/I1<4>/Q#3	VSS#263
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<3>/NM0	I0<5>/I1<3>/Q#6	WL#174	BL<44>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<3>/NM2	I0<5>/I1<3>/Q#6	I0<5>/I1<3>/QB#2	VSS#269
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<3>/NM1	BLB<44>#3	WL#180	I0<5>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<3>/NM3	I0<5>/I1<3>/QB#4	I0<5>/I1<3>/Q	VSS#276
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<2>/NM0	I0<5>/I1<2>/Q#4	WL#168	BL<41>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<2>/NM2	I0<5>/I1<2>/Q#4	I0<5>/I1<2>/QB	VSS#258
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<2>/NM1	BLB<41>#1	WL#162	I0<5>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<2>/NM3	I0<5>/I1<2>/QB#6	I0<5>/I1<2>/Q#3	VSS#251
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<1>/NM0	I0<5>/I1<1>/Q#6	WL#166	BL<42>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<1>/NM2	I0<5>/I1<1>/Q#6	I0<5>/I1<1>/QB#2	VSS#257
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<1>/NM1	BLB<42>#3	WL#172	I0<5>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<1>/NM3	I0<5>/I1<1>/QB#4	I0<5>/I1<1>/Q	VSS#264
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<0>/NM0	I0<5>/I1<0>/Q#6	WL#158	BL<40>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<0>/NM2	I0<5>/I1<0>/Q#6	I0<5>/I1<0>/QB#2	VSS#245
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<5>/I1<0>/NM1	BLB<40>#3	WL#164	I0<5>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<5>/I1<0>/NM3	I0<5>/I1<0>/QB#4	I0<5>/I1<0>/Q	VSS#252
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<7>/NM0	I0<4>/I1<7>/Q#4	WL#160	BL<39>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<7>/NM2	I0<4>/I1<7>/Q#4	I0<4>/I1<7>/QB	VSS#246
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<7>/NM1	BLB<39>#1	WL#154	I0<4>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<7>/NM3	I0<4>/I1<7>/QB#6	I0<4>/I1<7>/Q#3	VSS#239
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<6>/NM0	I0<4>/I1<6>/Q#4	WL#152	BL<37>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<6>/NM2	I0<4>/I1<6>/Q#4	I0<4>/I1<6>/QB	VSS#234
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<6>/NM1	BLB<37>#1	WL#146	I0<4>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<6>/NM3	I0<4>/I1<6>/QB#6	I0<4>/I1<6>/Q#3	VSS#227
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<5>/NM0	I0<4>/I1<5>/Q#6	WL#150	BL<38>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<5>/NM2	I0<4>/I1<5>/Q#6	I0<4>/I1<5>/QB#2	VSS#233
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<5>/NM1	BLB<38>#3	WL#156	I0<4>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<5>/NM3	I0<4>/I1<5>/QB#4	I0<4>/I1<5>/Q	VSS#240
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<4>/NM0	I0<4>/I1<4>/Q#4	WL#144	BL<35>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<4>/NM2	I0<4>/I1<4>/Q#4	I0<4>/I1<4>/QB	VSS#222
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<4>/NM1	BLB<35>#1	WL#138	I0<4>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<4>/NM3	I0<4>/I1<4>/QB#6	I0<4>/I1<4>/Q#3	VSS#215
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<3>/NM0	I0<4>/I1<3>/Q#6	WL#142	BL<36>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<3>/NM2	I0<4>/I1<3>/Q#6	I0<4>/I1<3>/QB#2	VSS#221
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<3>/NM1	BLB<36>#3	WL#148	I0<4>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<3>/NM3	I0<4>/I1<3>/QB#4	I0<4>/I1<3>/Q	VSS#228
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<2>/NM0	I0<4>/I1<2>/Q#4	WL#136	BL<33>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<2>/NM2	I0<4>/I1<2>/Q#4	I0<4>/I1<2>/QB	VSS#210
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<2>/NM1	BLB<33>#1	WL#130	I0<4>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<2>/NM3	I0<4>/I1<2>/QB#6	I0<4>/I1<2>/Q#3	VSS#203
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<1>/NM0	I0<4>/I1<1>/Q#6	WL#134	BL<34>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<1>/NM2	I0<4>/I1<1>/Q#6	I0<4>/I1<1>/QB#2	VSS#209
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<1>/NM1	BLB<34>#3	WL#140	I0<4>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<1>/NM3	I0<4>/I1<1>/QB#4	I0<4>/I1<1>/Q	VSS#216
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<0>/NM0	I0<4>/I1<0>/Q#6	WL#126	BL<32>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<0>/NM2	I0<4>/I1<0>/Q#6	I0<4>/I1<0>/QB#2	VSS#197
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<4>/I1<0>/NM1	BLB<32>#3	WL#132	I0<4>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<4>/I1<0>/NM3	I0<4>/I1<0>/QB#4	I0<4>/I1<0>/Q	VSS#204
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<7>/NM0	I0<3>/I1<7>/Q#4	WL#128	BL<31>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<7>/NM2	I0<3>/I1<7>/Q#4	I0<3>/I1<7>/QB	VSS#198
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<7>/NM1	BLB<31>#1	WL#122	I0<3>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<7>/NM3	I0<3>/I1<7>/QB#6	I0<3>/I1<7>/Q#3	VSS#191
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<6>/NM0	I0<3>/I1<6>/Q#4	WL#120	BL<29>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<6>/NM2	I0<3>/I1<6>/Q#4	I0<3>/I1<6>/QB	VSS#186
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<6>/NM1	BLB<29>#1	WL#114	I0<3>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<6>/NM3	I0<3>/I1<6>/QB#6	I0<3>/I1<6>/Q#3	VSS#179
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<5>/NM0	I0<3>/I1<5>/Q#6	WL#118	BL<30>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<5>/NM2	I0<3>/I1<5>/Q#6	I0<3>/I1<5>/QB#2	VSS#185
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<5>/NM1	BLB<30>#3	WL#124	I0<3>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<5>/NM3	I0<3>/I1<5>/QB#4	I0<3>/I1<5>/Q	VSS#192
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<4>/NM0	I0<3>/I1<4>/Q#4	WL#112	BL<27>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<4>/NM2	I0<3>/I1<4>/Q#4	I0<3>/I1<4>/QB	VSS#174
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<4>/NM1	BLB<27>#1	WL#106	I0<3>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<4>/NM3	I0<3>/I1<4>/QB#6	I0<3>/I1<4>/Q#3	VSS#167
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<3>/NM0	I0<3>/I1<3>/Q#6	WL#110	BL<28>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<3>/NM2	I0<3>/I1<3>/Q#6	I0<3>/I1<3>/QB#2	VSS#173
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<3>/NM1	BLB<28>#3	WL#116	I0<3>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<3>/NM3	I0<3>/I1<3>/QB#4	I0<3>/I1<3>/Q	VSS#180
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<2>/NM0	I0<3>/I1<2>/Q#4	WL#104	BL<25>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<2>/NM2	I0<3>/I1<2>/Q#4	I0<3>/I1<2>/QB	VSS#162
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<2>/NM1	BLB<25>#1	WL#98	I0<3>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<2>/NM3	I0<3>/I1<2>/QB#6	I0<3>/I1<2>/Q#3	VSS#155
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<1>/NM0	I0<3>/I1<1>/Q#6	WL#102	BL<26>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<1>/NM2	I0<3>/I1<1>/Q#6	I0<3>/I1<1>/QB#2	VSS#161
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<1>/NM1	BLB<26>#3	WL#108	I0<3>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<1>/NM3	I0<3>/I1<1>/QB#4	I0<3>/I1<1>/Q	VSS#168
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<0>/NM0	I0<3>/I1<0>/Q#6	WL#94	BL<24>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<0>/NM2	I0<3>/I1<0>/Q#6	I0<3>/I1<0>/QB#2	VSS#149
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<3>/I1<0>/NM1	BLB<24>#3	WL#100	I0<3>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<3>/I1<0>/NM3	I0<3>/I1<0>/QB#4	I0<3>/I1<0>/Q	VSS#156
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<7>/NM0	I0<2>/I1<7>/Q#4	WL#96	BL<23>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<7>/NM2	I0<2>/I1<7>/Q#4	I0<2>/I1<7>/QB	VSS#150
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<7>/NM1	BLB<23>#1	WL#90	I0<2>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<7>/NM3	I0<2>/I1<7>/QB#6	I0<2>/I1<7>/Q#3	VSS#143
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<6>/NM0	I0<2>/I1<6>/Q#4	WL#88	BL<21>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<6>/NM2	I0<2>/I1<6>/Q#4	I0<2>/I1<6>/QB	VSS#138
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<6>/NM1	BLB<21>#1	WL#82	I0<2>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<6>/NM3	I0<2>/I1<6>/QB#6	I0<2>/I1<6>/Q#3	VSS#131
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<5>/NM0	I0<2>/I1<5>/Q#6	WL#86	BL<22>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<5>/NM2	I0<2>/I1<5>/Q#6	I0<2>/I1<5>/QB#2	VSS#137
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<5>/NM1	BLB<22>#3	WL#92	I0<2>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<5>/NM3	I0<2>/I1<5>/QB#4	I0<2>/I1<5>/Q	VSS#144
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<4>/NM0	I0<2>/I1<4>/Q#4	WL#80	BL<19>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<4>/NM2	I0<2>/I1<4>/Q#4	I0<2>/I1<4>/QB	VSS#126
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<4>/NM1	BLB<19>#1	WL#74	I0<2>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<4>/NM3	I0<2>/I1<4>/QB#6	I0<2>/I1<4>/Q#3	VSS#119
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<3>/NM0	I0<2>/I1<3>/Q#6	WL#78	BL<20>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<3>/NM2	I0<2>/I1<3>/Q#6	I0<2>/I1<3>/QB#2	VSS#125
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<3>/NM1	BLB<20>#3	WL#84	I0<2>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<3>/NM3	I0<2>/I1<3>/QB#4	I0<2>/I1<3>/Q	VSS#132
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<2>/NM0	I0<2>/I1<2>/Q#4	WL#72	BL<17>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<2>/NM2	I0<2>/I1<2>/Q#4	I0<2>/I1<2>/QB	VSS#114
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<2>/NM1	BLB<17>#1	WL#66	I0<2>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<2>/NM3	I0<2>/I1<2>/QB#6	I0<2>/I1<2>/Q#3	VSS#107
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<1>/NM0	I0<2>/I1<1>/Q#6	WL#70	BL<18>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<1>/NM2	I0<2>/I1<1>/Q#6	I0<2>/I1<1>/QB#2	VSS#113
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<1>/NM1	BLB<18>#3	WL#76	I0<2>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<1>/NM3	I0<2>/I1<1>/QB#4	I0<2>/I1<1>/Q	VSS#120
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<0>/NM0	I0<2>/I1<0>/Q#6	WL#62	BL<16>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<0>/NM2	I0<2>/I1<0>/Q#6	I0<2>/I1<0>/QB#2	VSS#101
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<2>/I1<0>/NM1	BLB<16>#3	WL#68	I0<2>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<2>/I1<0>/NM3	I0<2>/I1<0>/QB#4	I0<2>/I1<0>/Q	VSS#108
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<7>/NM0	I0<1>/I1<7>/Q#4	WL#64	BL<15>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<7>/NM2	I0<1>/I1<7>/Q#4	I0<1>/I1<7>/QB	VSS#102
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<7>/NM1	BLB<15>#1	WL#58	I0<1>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<7>/NM3	I0<1>/I1<7>/QB#6	I0<1>/I1<7>/Q#3	VSS#95
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<6>/NM0	I0<1>/I1<6>/Q#4	WL#56	BL<13>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<6>/NM2	I0<1>/I1<6>/Q#4	I0<1>/I1<6>/QB	VSS#90	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<6>/NM1	BLB<13>#1	WL#50	I0<1>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<6>/NM3	I0<1>/I1<6>/QB#6	I0<1>/I1<6>/Q#3	VSS#83
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<5>/NM0	I0<1>/I1<5>/Q#6	WL#54	BL<14>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<5>/NM2	I0<1>/I1<5>/Q#6	I0<1>/I1<5>/QB#2	VSS#89
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<5>/NM1	BLB<14>#3	WL#60	I0<1>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<5>/NM3	I0<1>/I1<5>/QB#4	I0<1>/I1<5>/Q	VSS#96	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<4>/NM0	I0<1>/I1<4>/Q#4	WL#48	BL<11>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<4>/NM2	I0<1>/I1<4>/Q#4	I0<1>/I1<4>/QB	VSS#78	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<4>/NM1	BLB<11>#1	WL#42	I0<1>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<4>/NM3	I0<1>/I1<4>/QB#6	I0<1>/I1<4>/Q#3	VSS#71
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<3>/NM0	I0<1>/I1<3>/Q#6	WL#46	BL<12>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<3>/NM2	I0<1>/I1<3>/Q#6	I0<1>/I1<3>/QB#2	VSS#77
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<3>/NM1	BLB<12>#3	WL#52	I0<1>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<3>/NM3	I0<1>/I1<3>/QB#4	I0<1>/I1<3>/Q	VSS#84	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<2>/NM0	I0<1>/I1<2>/Q#4	WL#40	BL<9>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<2>/NM2	I0<1>/I1<2>/Q#4	I0<1>/I1<2>/QB	VSS#66	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<2>/NM1	BLB<9>#1	WL#34	I0<1>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<2>/NM3	I0<1>/I1<2>/QB#6	I0<1>/I1<2>/Q#3	VSS#59
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<1>/NM0	I0<1>/I1<1>/Q#6	WL#38	BL<10>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<1>/NM2	I0<1>/I1<1>/Q#6	I0<1>/I1<1>/QB#2	VSS#65
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<1>/NM1	BLB<10>#3	WL#44	I0<1>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<1>/NM3	I0<1>/I1<1>/QB#4	I0<1>/I1<1>/Q	VSS#72	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<0>/NM0	I0<1>/I1<0>/Q#6	WL#30	BL<8>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<0>/NM2	I0<1>/I1<0>/Q#6	I0<1>/I1<0>/QB#2	VSS#53
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<1>/I1<0>/NM1	BLB<8>#3	WL#36	I0<1>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<1>/I1<0>/NM3	I0<1>/I1<0>/QB#4	I0<1>/I1<0>/Q	VSS#60	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<7>/NM0	I0<0>/I1<7>/Q#4	WL#32	BL<7>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<7>/NM2	I0<0>/I1<7>/Q#4	I0<0>/I1<7>/QB	VSS#54	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<7>/NM1	BLB<7>#1	WL#26	I0<0>/I1<7>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<7>/NM3	I0<0>/I1<7>/QB#6	I0<0>/I1<7>/Q#3	VSS#47
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<6>/NM0	I0<0>/I1<6>/Q#4	WL#24	BL<5>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<6>/NM2	I0<0>/I1<6>/Q#4	I0<0>/I1<6>/QB	VSS#42	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<6>/NM1	BLB<5>#1	WL#18	I0<0>/I1<6>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<6>/NM3	I0<0>/I1<6>/QB#6	I0<0>/I1<6>/Q#3	VSS#35
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<5>/NM0	I0<0>/I1<5>/Q#6	WL#22	BL<6>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<5>/NM2	I0<0>/I1<5>/Q#6	I0<0>/I1<5>/QB#2	VSS#41
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<5>/NM1	BLB<6>#3	WL#28	I0<0>/I1<5>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<5>/NM3	I0<0>/I1<5>/QB#4	I0<0>/I1<5>/Q	VSS#48	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<4>/NM0	I0<0>/I1<4>/Q#4	WL#16	BL<3>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<4>/NM2	I0<0>/I1<4>/Q#4	I0<0>/I1<4>/QB	VSS#30	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<4>/NM1	BLB<3>#1	WL#10	I0<0>/I1<4>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<4>/NM3	I0<0>/I1<4>/QB#6	I0<0>/I1<4>/Q#3	VSS#23
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<3>/NM0	I0<0>/I1<3>/Q#6	WL#14	BL<4>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<3>/NM2	I0<0>/I1<3>/Q#6	I0<0>/I1<3>/QB#2	VSS#29
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<3>/NM1	BLB<4>#3	WL#20	I0<0>/I1<3>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<3>/NM3	I0<0>/I1<3>/QB#4	I0<0>/I1<3>/Q	VSS#36	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<2>/NM0	I0<0>/I1<2>/Q#4	WL#8	BL<1>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<2>/NM2	I0<0>/I1<2>/Q#4	I0<0>/I1<2>/QB	VSS#18	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<2>/NM1	BLB<1>#1	WL#3	I0<0>/I1<2>/QB#6	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<2>/NM3	I0<0>/I1<2>/QB#6	I0<0>/I1<2>/Q#3	VSS#11
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<1>/NM0	I0<0>/I1<1>/Q#6	WL#6	BL<2>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<1>/NM2	I0<0>/I1<1>/Q#6	I0<0>/I1<1>/QB#2	VSS#17
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<1>/NM1	BLB<2>#3	WL#12	I0<0>/I1<1>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<1>/NM3	I0<0>/I1<1>/QB#4	I0<0>/I1<1>/Q	VSS#24	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<0>/NM0	I0<0>/I1<0>/Q#6	WL#1	BL<0>#1	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<0>/NM2	I0<0>/I1<0>/Q#6	I0<0>/I1<0>/QB#2	VSS#6
+ VSS#4	nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<0>/I1<0>/NM1	BLB<0>#3	WL#5	I0<0>/I1<0>/QB#4	VSS#4
+ nmos1v	L=4.5e-08	W=1.2e-07
+ AD=2.75e-14	AS=2.75e-14	PD=6.8e-07	PS=6.8e-07
MI0<0>/I1<0>/NM3	I0<0>/I1<0>/QB#4	I0<0>/I1<0>/Q	VSS#12	VSS#4
+ nmos1v	L=4.5e-08	W=2.3e-07
+ AD=3.52e-14	AS=3.52e-14	PD=7.9e-07	PS=7.9e-07
MI0<7>/I1<7>/PM0	I0<7>/I1<7>/Q#5	I0<7>/I1<7>/QB#2	VDD#566
+ VDD#565	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<7>/PM1	I0<7>/I1<7>/QB#4	I0<7>/I1<7>/Q#2	VDD#563
+ VDD#565	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<6>/PM0	I0<7>/I1<6>/Q#5	I0<7>/I1<6>/QB#2	VDD#554
+ VDD#553	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<6>/PM1	I0<7>/I1<6>/QB#4	I0<7>/I1<6>/Q#2	VDD#551
+ VDD#553	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<5>/PM0	I0<7>/I1<5>/Q#4	I0<7>/I1<5>/QB	VDD#557
+ VDD#559	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<5>/PM1	I0<7>/I1<5>/QB#5	I0<7>/I1<5>/Q#2	VDD#560
+ VDD#559	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<4>/PM0	I0<7>/I1<4>/Q#5	I0<7>/I1<4>/QB#2	VDD#536
+ VDD#535	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<4>/PM1	I0<7>/I1<4>/QB#4	I0<7>/I1<4>/Q#2	VDD#533
+ VDD#535	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<3>/PM0	I0<7>/I1<3>/Q#4	I0<7>/I1<3>/QB	VDD#542
+ VDD#544	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<3>/PM1	I0<7>/I1<3>/QB#5	I0<7>/I1<3>/Q#2	VDD#545
+ VDD#544	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<2>/PM0	I0<7>/I1<2>/Q#5	I0<7>/I1<2>/QB#2	VDD#518
+ VDD#517	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<2>/PM1	I0<7>/I1<2>/QB#4	I0<7>/I1<2>/Q#2	VDD#515
+ VDD#517	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<1>/PM0	I0<7>/I1<1>/Q#4	I0<7>/I1<1>/QB	VDD#524
+ VDD#526	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<1>/PM1	I0<7>/I1<1>/QB#5	I0<7>/I1<1>/Q#2	VDD#527
+ VDD#526	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<0>/PM0	I0<7>/I1<0>/Q#4	I0<7>/I1<0>/QB	VDD#506
+ VDD#508	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<7>/I1<0>/PM1	I0<7>/I1<0>/QB#5	I0<7>/I1<0>/Q#2	VDD#509
+ VDD#508	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<7>/PM0	I0<6>/I1<7>/Q#5	I0<6>/I1<7>/QB#2	VDD#500
+ VDD#499	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<7>/PM1	I0<6>/I1<7>/QB#4	I0<6>/I1<7>/Q#2	VDD#497
+ VDD#499	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<6>/PM0	I0<6>/I1<6>/Q#5	I0<6>/I1<6>/QB#2	VDD#482
+ VDD#481	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<6>/PM1	I0<6>/I1<6>/QB#4	I0<6>/I1<6>/Q#2	VDD#479
+ VDD#481	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<5>/PM0	I0<6>/I1<5>/Q#4	I0<6>/I1<5>/QB	VDD#488
+ VDD#490	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<5>/PM1	I0<6>/I1<5>/QB#5	I0<6>/I1<5>/Q#2	VDD#491
+ VDD#490	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<4>/PM0	I0<6>/I1<4>/Q#5	I0<6>/I1<4>/QB#2	VDD#464
+ VDD#463	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<4>/PM1	I0<6>/I1<4>/QB#4	I0<6>/I1<4>/Q#2	VDD#461
+ VDD#463	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<3>/PM0	I0<6>/I1<3>/Q#4	I0<6>/I1<3>/QB	VDD#470
+ VDD#472	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<3>/PM1	I0<6>/I1<3>/QB#5	I0<6>/I1<3>/Q#2	VDD#473
+ VDD#472	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<2>/PM0	I0<6>/I1<2>/Q#5	I0<6>/I1<2>/QB#2	VDD#446
+ VDD#445	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<2>/PM1	I0<6>/I1<2>/QB#4	I0<6>/I1<2>/Q#2	VDD#443
+ VDD#445	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<1>/PM0	I0<6>/I1<1>/Q#4	I0<6>/I1<1>/QB	VDD#452
+ VDD#454	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<1>/PM1	I0<6>/I1<1>/QB#5	I0<6>/I1<1>/Q#2	VDD#455
+ VDD#454	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<0>/PM0	I0<6>/I1<0>/Q#4	I0<6>/I1<0>/QB	VDD#434
+ VDD#436	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<6>/I1<0>/PM1	I0<6>/I1<0>/QB#5	I0<6>/I1<0>/Q#2	VDD#437
+ VDD#436	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<7>/PM0	I0<5>/I1<7>/Q#5	I0<5>/I1<7>/QB#2	VDD#428
+ VDD#427	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<7>/PM1	I0<5>/I1<7>/QB#4	I0<5>/I1<7>/Q#2	VDD#425
+ VDD#427	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<6>/PM0	I0<5>/I1<6>/Q#5	I0<5>/I1<6>/QB#2	VDD#410
+ VDD#409	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<6>/PM1	I0<5>/I1<6>/QB#4	I0<5>/I1<6>/Q#2	VDD#407
+ VDD#409	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<5>/PM0	I0<5>/I1<5>/Q#4	I0<5>/I1<5>/QB	VDD#416
+ VDD#418	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<5>/PM1	I0<5>/I1<5>/QB#5	I0<5>/I1<5>/Q#2	VDD#419
+ VDD#418	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<4>/PM0	I0<5>/I1<4>/Q#5	I0<5>/I1<4>/QB#2	VDD#392
+ VDD#391	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<4>/PM1	I0<5>/I1<4>/QB#4	I0<5>/I1<4>/Q#2	VDD#389
+ VDD#391	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<3>/PM0	I0<5>/I1<3>/Q#4	I0<5>/I1<3>/QB	VDD#398
+ VDD#400	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<3>/PM1	I0<5>/I1<3>/QB#5	I0<5>/I1<3>/Q#2	VDD#401
+ VDD#400	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<2>/PM0	I0<5>/I1<2>/Q#5	I0<5>/I1<2>/QB#2	VDD#374
+ VDD#373	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<2>/PM1	I0<5>/I1<2>/QB#4	I0<5>/I1<2>/Q#2	VDD#371
+ VDD#373	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<1>/PM0	I0<5>/I1<1>/Q#4	I0<5>/I1<1>/QB	VDD#380
+ VDD#382	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<1>/PM1	I0<5>/I1<1>/QB#5	I0<5>/I1<1>/Q#2	VDD#383
+ VDD#382	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<0>/PM0	I0<5>/I1<0>/Q#4	I0<5>/I1<0>/QB	VDD#362
+ VDD#364	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<5>/I1<0>/PM1	I0<5>/I1<0>/QB#5	I0<5>/I1<0>/Q#2	VDD#365
+ VDD#364	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<7>/PM0	I0<4>/I1<7>/Q#5	I0<4>/I1<7>/QB#2	VDD#356
+ VDD#355	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<7>/PM1	I0<4>/I1<7>/QB#4	I0<4>/I1<7>/Q#2	VDD#353
+ VDD#355	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<6>/PM0	I0<4>/I1<6>/Q#5	I0<4>/I1<6>/QB#2	VDD#338
+ VDD#337	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<6>/PM1	I0<4>/I1<6>/QB#4	I0<4>/I1<6>/Q#2	VDD#335
+ VDD#337	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<5>/PM0	I0<4>/I1<5>/Q#4	I0<4>/I1<5>/QB	VDD#344
+ VDD#346	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<5>/PM1	I0<4>/I1<5>/QB#5	I0<4>/I1<5>/Q#2	VDD#347
+ VDD#346	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<4>/PM0	I0<4>/I1<4>/Q#5	I0<4>/I1<4>/QB#2	VDD#320
+ VDD#319	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<4>/PM1	I0<4>/I1<4>/QB#4	I0<4>/I1<4>/Q#2	VDD#317
+ VDD#319	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<3>/PM0	I0<4>/I1<3>/Q#4	I0<4>/I1<3>/QB	VDD#326
+ VDD#328	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<3>/PM1	I0<4>/I1<3>/QB#5	I0<4>/I1<3>/Q#2	VDD#329
+ VDD#328	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<2>/PM0	I0<4>/I1<2>/Q#5	I0<4>/I1<2>/QB#2	VDD#302
+ VDD#301	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<2>/PM1	I0<4>/I1<2>/QB#4	I0<4>/I1<2>/Q#2	VDD#299
+ VDD#301	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<1>/PM0	I0<4>/I1<1>/Q#4	I0<4>/I1<1>/QB	VDD#308
+ VDD#310	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<1>/PM1	I0<4>/I1<1>/QB#5	I0<4>/I1<1>/Q#2	VDD#311
+ VDD#310	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<0>/PM0	I0<4>/I1<0>/Q#4	I0<4>/I1<0>/QB	VDD#290
+ VDD#292	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<4>/I1<0>/PM1	I0<4>/I1<0>/QB#5	I0<4>/I1<0>/Q#2	VDD#293
+ VDD#292	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<7>/PM0	I0<3>/I1<7>/Q#5	I0<3>/I1<7>/QB#2	VDD#284
+ VDD#283	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<7>/PM1	I0<3>/I1<7>/QB#4	I0<3>/I1<7>/Q#2	VDD#281
+ VDD#283	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<6>/PM0	I0<3>/I1<6>/Q#5	I0<3>/I1<6>/QB#2	VDD#266
+ VDD#265	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<6>/PM1	I0<3>/I1<6>/QB#4	I0<3>/I1<6>/Q#2	VDD#263
+ VDD#265	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<5>/PM0	I0<3>/I1<5>/Q#4	I0<3>/I1<5>/QB	VDD#272
+ VDD#274	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<5>/PM1	I0<3>/I1<5>/QB#5	I0<3>/I1<5>/Q#2	VDD#275
+ VDD#274	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<4>/PM0	I0<3>/I1<4>/Q#5	I0<3>/I1<4>/QB#2	VDD#248
+ VDD#247	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<4>/PM1	I0<3>/I1<4>/QB#4	I0<3>/I1<4>/Q#2	VDD#245
+ VDD#247	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<3>/PM0	I0<3>/I1<3>/Q#4	I0<3>/I1<3>/QB	VDD#254
+ VDD#256	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<3>/PM1	I0<3>/I1<3>/QB#5	I0<3>/I1<3>/Q#2	VDD#257
+ VDD#256	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<2>/PM0	I0<3>/I1<2>/Q#5	I0<3>/I1<2>/QB#2	VDD#230
+ VDD#229	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<2>/PM1	I0<3>/I1<2>/QB#4	I0<3>/I1<2>/Q#2	VDD#227
+ VDD#229	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<1>/PM0	I0<3>/I1<1>/Q#4	I0<3>/I1<1>/QB	VDD#236
+ VDD#238	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<1>/PM1	I0<3>/I1<1>/QB#5	I0<3>/I1<1>/Q#2	VDD#239
+ VDD#238	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<0>/PM0	I0<3>/I1<0>/Q#4	I0<3>/I1<0>/QB	VDD#218
+ VDD#220	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<3>/I1<0>/PM1	I0<3>/I1<0>/QB#5	I0<3>/I1<0>/Q#2	VDD#221
+ VDD#220	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<7>/PM0	I0<2>/I1<7>/Q#5	I0<2>/I1<7>/QB#2	VDD#212
+ VDD#211	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<7>/PM1	I0<2>/I1<7>/QB#4	I0<2>/I1<7>/Q#2	VDD#209
+ VDD#211	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<6>/PM0	I0<2>/I1<6>/Q#5	I0<2>/I1<6>/QB#2	VDD#194
+ VDD#193	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<6>/PM1	I0<2>/I1<6>/QB#4	I0<2>/I1<6>/Q#2	VDD#191
+ VDD#193	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<5>/PM0	I0<2>/I1<5>/Q#4	I0<2>/I1<5>/QB	VDD#200
+ VDD#202	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<5>/PM1	I0<2>/I1<5>/QB#5	I0<2>/I1<5>/Q#2	VDD#203
+ VDD#202	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<4>/PM0	I0<2>/I1<4>/Q#5	I0<2>/I1<4>/QB#2	VDD#176
+ VDD#175	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<4>/PM1	I0<2>/I1<4>/QB#4	I0<2>/I1<4>/Q#2	VDD#173
+ VDD#175	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<3>/PM0	I0<2>/I1<3>/Q#4	I0<2>/I1<3>/QB	VDD#182
+ VDD#184	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<3>/PM1	I0<2>/I1<3>/QB#5	I0<2>/I1<3>/Q#2	VDD#185
+ VDD#184	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<2>/PM0	I0<2>/I1<2>/Q#5	I0<2>/I1<2>/QB#2	VDD#158
+ VDD#157	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<2>/PM1	I0<2>/I1<2>/QB#4	I0<2>/I1<2>/Q#2	VDD#155
+ VDD#157	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<1>/PM0	I0<2>/I1<1>/Q#4	I0<2>/I1<1>/QB	VDD#164
+ VDD#166	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<1>/PM1	I0<2>/I1<1>/QB#5	I0<2>/I1<1>/Q#2	VDD#167
+ VDD#166	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<0>/PM0	I0<2>/I1<0>/Q#4	I0<2>/I1<0>/QB	VDD#146
+ VDD#148	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<2>/I1<0>/PM1	I0<2>/I1<0>/QB#5	I0<2>/I1<0>/Q#2	VDD#149
+ VDD#148	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<7>/PM0	I0<1>/I1<7>/Q#5	I0<1>/I1<7>/QB#2	VDD#140
+ VDD#139	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<7>/PM1	I0<1>/I1<7>/QB#4	I0<1>/I1<7>/Q#2	VDD#137
+ VDD#139	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<6>/PM0	I0<1>/I1<6>/Q#5	I0<1>/I1<6>/QB#2	VDD#122
+ VDD#121	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<6>/PM1	I0<1>/I1<6>/QB#4	I0<1>/I1<6>/Q#2	VDD#119
+ VDD#121	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<5>/PM0	I0<1>/I1<5>/Q#4	I0<1>/I1<5>/QB	VDD#128
+ VDD#130	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<5>/PM1	I0<1>/I1<5>/QB#5	I0<1>/I1<5>/Q#2	VDD#131
+ VDD#130	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<4>/PM0	I0<1>/I1<4>/Q#5	I0<1>/I1<4>/QB#2	VDD#104
+ VDD#103	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<4>/PM1	I0<1>/I1<4>/QB#4	I0<1>/I1<4>/Q#2	VDD#101
+ VDD#103	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<3>/PM0	I0<1>/I1<3>/Q#4	I0<1>/I1<3>/QB	VDD#110
+ VDD#112	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<3>/PM1	I0<1>/I1<3>/QB#5	I0<1>/I1<3>/Q#2	VDD#113
+ VDD#112	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<2>/PM0	I0<1>/I1<2>/Q#5	I0<1>/I1<2>/QB#2	VDD#86
+ VDD#85	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<2>/PM1	I0<1>/I1<2>/QB#4	I0<1>/I1<2>/Q#2	VDD#83
+ VDD#85	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<1>/PM0	I0<1>/I1<1>/Q#4	I0<1>/I1<1>/QB	VDD#92	VDD#94
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<1>/PM1	I0<1>/I1<1>/QB#5	I0<1>/I1<1>/Q#2	VDD#95
+ VDD#94	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<0>/PM0	I0<1>/I1<0>/Q#4	I0<1>/I1<0>/QB	VDD#74	VDD#76
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<1>/I1<0>/PM1	I0<1>/I1<0>/QB#5	I0<1>/I1<0>/Q#2	VDD#77
+ VDD#76	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<7>/PM0	I0<0>/I1<7>/Q#5	I0<0>/I1<7>/QB#2	VDD#68
+ VDD#67	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<7>/PM1	I0<0>/I1<7>/QB#4	I0<0>/I1<7>/Q#2	VDD#65
+ VDD#67	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<6>/PM0	I0<0>/I1<6>/Q#5	I0<0>/I1<6>/QB#2	VDD#50
+ VDD#49	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<6>/PM1	I0<0>/I1<6>/QB#4	I0<0>/I1<6>/Q#2	VDD#47
+ VDD#49	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<5>/PM0	I0<0>/I1<5>/Q#4	I0<0>/I1<5>/QB	VDD#56	VDD#58
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<5>/PM1	I0<0>/I1<5>/QB#5	I0<0>/I1<5>/Q#2	VDD#59
+ VDD#58	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<4>/PM0	I0<0>/I1<4>/Q#5	I0<0>/I1<4>/QB#2	VDD#32
+ VDD#31	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<4>/PM1	I0<0>/I1<4>/QB#4	I0<0>/I1<4>/Q#2	VDD#29
+ VDD#31	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<3>/PM0	I0<0>/I1<3>/Q#4	I0<0>/I1<3>/QB	VDD#38	VDD#40
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<3>/PM1	I0<0>/I1<3>/QB#5	I0<0>/I1<3>/Q#2	VDD#41
+ VDD#40	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<2>/PM0	I0<0>/I1<2>/Q#5	I0<0>/I1<2>/QB#2	VDD#14
+ VDD#13	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<2>/PM1	I0<0>/I1<2>/QB#4	I0<0>/I1<2>/Q#2	VDD#11
+ VDD#13	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<1>/PM0	I0<0>/I1<1>/Q#4	I0<0>/I1<1>/QB	VDD#20	VDD#22
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<1>/PM1	I0<0>/I1<1>/QB#5	I0<0>/I1<1>/Q#2	VDD#23
+ VDD#22	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<0>/PM0	I0<0>/I1<0>/Q#4	I0<0>/I1<0>/QB	VDD#2	VDD#4
+ pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
MI0<0>/I1<0>/PM1	I0<0>/I1<0>/QB#5	I0<0>/I1<0>/Q#2	VDD#5
+ VDD#4	pmos1v	L=4.5e-08	W=1.2e-07
+ AD=1.68e-14	AS=1.68e-14	PD=5.2e-07	PS=5.2e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	WL#1	WL#2	  104.7064	$poly_conn
Rl2	I0<0>/I1<0>/QB	I0<0>/I1<0>/QB#2	   56.4103	$poly_conn
Rl3	I0<0>/I1<0>/QB	I0<0>/I1<0>/QB#3	   90.3330	$poly_conn
Rl4	I0<0>/I1<0>/Q	I0<0>/I1<0>/Q#2	   56.4103	$poly_conn
Rl5	I0<0>/I1<0>/Q#2	I0<0>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl6	WL#3	WL#4	   59.7064	$poly_conn
Rl7	WL#4	WL#5	   59.7064	$poly_conn
Rl8	I0<0>/I1<2>/Q	I0<0>/I1<2>/Q#2	   90.3330	$poly_conn
Rl9	I0<0>/I1<2>/Q#2	I0<0>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl10	I0<0>/I1<2>/QB	I0<0>/I1<2>/QB#2	   56.4103	$poly_conn
Rl11	I0<0>/I1<2>/QB#2	I0<0>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl12	WL#6	WL#7	   59.7064	$poly_conn
Rl13	WL#7	WL#8	   59.7064	$poly_conn
Rl14	I0<0>/I1<1>/QB	I0<0>/I1<1>/QB#2	   56.4103	$poly_conn
Rl15	I0<0>/I1<1>/QB	I0<0>/I1<1>/QB#3	   90.3330	$poly_conn
Rl16	I0<0>/I1<1>/Q	I0<0>/I1<1>/Q#2	   56.4103	$poly_conn
Rl17	I0<0>/I1<1>/Q#2	I0<0>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl18	WL#10	WL#11	   59.7064	$poly_conn
Rl19	WL#11	WL#12	   59.7064	$poly_conn
Rl20	I0<0>/I1<4>/Q	I0<0>/I1<4>/Q#2	   90.3330	$poly_conn
Rl21	I0<0>/I1<4>/Q#2	I0<0>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl22	I0<0>/I1<4>/QB	I0<0>/I1<4>/QB#2	   56.4103	$poly_conn
Rl23	I0<0>/I1<4>/QB#2	I0<0>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl24	WL#14	WL#15	   59.7064	$poly_conn
Rl25	WL#15	WL#16	   59.7064	$poly_conn
Rl26	I0<0>/I1<3>/QB	I0<0>/I1<3>/QB#2	   56.4103	$poly_conn
Rl27	I0<0>/I1<3>/QB	I0<0>/I1<3>/QB#3	   90.3330	$poly_conn
Rl28	I0<0>/I1<3>/Q	I0<0>/I1<3>/Q#2	   56.4103	$poly_conn
Rl29	I0<0>/I1<3>/Q#2	I0<0>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl30	WL#18	WL#19	   59.7064	$poly_conn
Rl31	WL#19	WL#20	   59.7064	$poly_conn
Rl32	I0<0>/I1<6>/Q	I0<0>/I1<6>/Q#2	   90.3330	$poly_conn
Rl33	I0<0>/I1<6>/Q#2	I0<0>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl34	I0<0>/I1<6>/QB	I0<0>/I1<6>/QB#2	   56.4103	$poly_conn
Rl35	I0<0>/I1<6>/QB#2	I0<0>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl36	WL#22	WL#23	   59.7064	$poly_conn
Rl37	WL#23	WL#24	   59.7064	$poly_conn
Rl38	I0<0>/I1<5>/QB	I0<0>/I1<5>/QB#2	   56.4103	$poly_conn
Rl39	I0<0>/I1<5>/QB	I0<0>/I1<5>/QB#3	   90.3330	$poly_conn
Rl40	I0<0>/I1<5>/Q	I0<0>/I1<5>/Q#2	   56.4103	$poly_conn
Rl41	I0<0>/I1<5>/Q#2	I0<0>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl42	WL#26	WL#27	   59.7064	$poly_conn
Rl43	WL#27	WL#28	   59.7064	$poly_conn
Rl44	I0<0>/I1<7>/Q	I0<0>/I1<7>/Q#2	   90.3330	$poly_conn
Rl45	I0<0>/I1<7>/Q#2	I0<0>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl46	I0<0>/I1<7>/QB	I0<0>/I1<7>/QB#2	   56.4103	$poly_conn
Rl47	I0<0>/I1<7>/QB#2	I0<0>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl48	WL#30	WL#31	   59.7064	$poly_conn
Rl49	WL#31	WL#32	   59.7064	$poly_conn
Rl50	I0<1>/I1<0>/QB	I0<1>/I1<0>/QB#2	   56.4103	$poly_conn
Rl51	I0<1>/I1<0>/QB	I0<1>/I1<0>/QB#3	   90.3330	$poly_conn
Rl52	I0<1>/I1<0>/Q	I0<1>/I1<0>/Q#2	   56.4103	$poly_conn
Rl53	I0<1>/I1<0>/Q#2	I0<1>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl54	WL#34	WL#35	   59.7064	$poly_conn
Rl55	WL#35	WL#36	   59.7064	$poly_conn
Rl56	I0<1>/I1<2>/Q	I0<1>/I1<2>/Q#2	   90.3330	$poly_conn
Rl57	I0<1>/I1<2>/Q#2	I0<1>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl58	I0<1>/I1<2>/QB	I0<1>/I1<2>/QB#2	   56.4103	$poly_conn
Rl59	I0<1>/I1<2>/QB#2	I0<1>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl60	WL#38	WL#39	   59.7064	$poly_conn
Rl61	WL#39	WL#40	   59.7064	$poly_conn
Rl62	I0<1>/I1<1>/QB	I0<1>/I1<1>/QB#2	   56.4103	$poly_conn
Rl63	I0<1>/I1<1>/QB	I0<1>/I1<1>/QB#3	   90.3330	$poly_conn
Rl64	I0<1>/I1<1>/Q	I0<1>/I1<1>/Q#2	   56.4103	$poly_conn
Rl65	I0<1>/I1<1>/Q#2	I0<1>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl66	WL#42	WL#43	   59.7064	$poly_conn
Rl67	WL#43	WL#44	   59.7064	$poly_conn
Rl68	I0<1>/I1<4>/Q	I0<1>/I1<4>/Q#2	   90.3330	$poly_conn
Rl69	I0<1>/I1<4>/Q#2	I0<1>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl70	I0<1>/I1<4>/QB	I0<1>/I1<4>/QB#2	   56.4103	$poly_conn
Rl71	I0<1>/I1<4>/QB#2	I0<1>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl72	WL#46	WL#47	   59.7064	$poly_conn
Rl73	WL#47	WL#48	   59.7064	$poly_conn
Rl74	I0<1>/I1<3>/QB	I0<1>/I1<3>/QB#2	   56.4103	$poly_conn
Rl75	I0<1>/I1<3>/QB	I0<1>/I1<3>/QB#3	   90.3330	$poly_conn
Rl76	I0<1>/I1<3>/Q	I0<1>/I1<3>/Q#2	   56.4103	$poly_conn
Rl77	I0<1>/I1<3>/Q#2	I0<1>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl78	WL#50	WL#51	   59.7064	$poly_conn
Rl79	WL#51	WL#52	   59.7064	$poly_conn
Rl80	I0<1>/I1<6>/Q	I0<1>/I1<6>/Q#2	   90.3330	$poly_conn
Rl81	I0<1>/I1<6>/Q#2	I0<1>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl82	I0<1>/I1<6>/QB	I0<1>/I1<6>/QB#2	   56.4103	$poly_conn
Rl83	I0<1>/I1<6>/QB#2	I0<1>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl84	WL#54	WL#55	   59.7064	$poly_conn
Rl85	WL#55	WL#56	   59.7064	$poly_conn
Rl86	I0<1>/I1<5>/QB	I0<1>/I1<5>/QB#2	   56.4103	$poly_conn
Rl87	I0<1>/I1<5>/QB	I0<1>/I1<5>/QB#3	   90.3330	$poly_conn
Rl88	I0<1>/I1<5>/Q	I0<1>/I1<5>/Q#2	   56.4103	$poly_conn
Rl89	I0<1>/I1<5>/Q#2	I0<1>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl90	WL#58	WL#59	   59.7064	$poly_conn
Rl91	WL#59	WL#60	   59.7064	$poly_conn
Rl92	I0<1>/I1<7>/Q	I0<1>/I1<7>/Q#2	   90.3330	$poly_conn
Rl93	I0<1>/I1<7>/Q#2	I0<1>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl94	I0<1>/I1<7>/QB	I0<1>/I1<7>/QB#2	   56.4103	$poly_conn
Rl95	I0<1>/I1<7>/QB#2	I0<1>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl96	WL#62	WL#63	   59.7064	$poly_conn
Rl97	WL#63	WL#64	   59.7064	$poly_conn
Rl98	I0<2>/I1<0>/QB	I0<2>/I1<0>/QB#2	   56.4103	$poly_conn
Rl99	I0<2>/I1<0>/QB	I0<2>/I1<0>/QB#3	   90.3330	$poly_conn
Rl100	I0<2>/I1<0>/Q	I0<2>/I1<0>/Q#2	   56.4103	$poly_conn
Rl101	I0<2>/I1<0>/Q#2	I0<2>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl102	WL#66	WL#67	   59.7064	$poly_conn
Rl103	WL#67	WL#68	   59.7064	$poly_conn
Rl104	I0<2>/I1<2>/Q	I0<2>/I1<2>/Q#2	   90.3330	$poly_conn
Rl105	I0<2>/I1<2>/Q#2	I0<2>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl106	I0<2>/I1<2>/QB	I0<2>/I1<2>/QB#2	   56.4103	$poly_conn
Rl107	I0<2>/I1<2>/QB#2	I0<2>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl108	WL#70	WL#71	   59.7064	$poly_conn
Rl109	WL#71	WL#72	   59.7064	$poly_conn
Rl110	I0<2>/I1<1>/QB	I0<2>/I1<1>/QB#2	   56.4103	$poly_conn
Rl111	I0<2>/I1<1>/QB	I0<2>/I1<1>/QB#3	   90.3330	$poly_conn
Rl112	I0<2>/I1<1>/Q	I0<2>/I1<1>/Q#2	   56.4103	$poly_conn
Rl113	I0<2>/I1<1>/Q#2	I0<2>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl114	WL#74	WL#75	   59.7064	$poly_conn
Rl115	WL#75	WL#76	   59.7064	$poly_conn
Rl116	I0<2>/I1<4>/Q	I0<2>/I1<4>/Q#2	   90.3330	$poly_conn
Rl117	I0<2>/I1<4>/Q#2	I0<2>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl118	I0<2>/I1<4>/QB	I0<2>/I1<4>/QB#2	   56.4103	$poly_conn
Rl119	I0<2>/I1<4>/QB#2	I0<2>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl120	WL#78	WL#79	   59.7064	$poly_conn
Rl121	WL#79	WL#80	   59.7064	$poly_conn
Rl122	I0<2>/I1<3>/QB	I0<2>/I1<3>/QB#2	   56.4103	$poly_conn
Rl123	I0<2>/I1<3>/QB	I0<2>/I1<3>/QB#3	   90.3330	$poly_conn
Rl124	I0<2>/I1<3>/Q	I0<2>/I1<3>/Q#2	   56.4103	$poly_conn
Rl125	I0<2>/I1<3>/Q#2	I0<2>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl126	WL#82	WL#83	   59.7064	$poly_conn
Rl127	WL#83	WL#84	   59.7064	$poly_conn
Rl128	I0<2>/I1<6>/Q	I0<2>/I1<6>/Q#2	   90.3330	$poly_conn
Rl129	I0<2>/I1<6>/Q#2	I0<2>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl130	I0<2>/I1<6>/QB	I0<2>/I1<6>/QB#2	   56.4103	$poly_conn
Rl131	I0<2>/I1<6>/QB#2	I0<2>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl132	WL#86	WL#87	   59.7064	$poly_conn
Rl133	WL#87	WL#88	   59.7064	$poly_conn
Rl134	I0<2>/I1<5>/QB	I0<2>/I1<5>/QB#2	   56.4103	$poly_conn
Rl135	I0<2>/I1<5>/QB	I0<2>/I1<5>/QB#3	   90.3330	$poly_conn
Rl136	I0<2>/I1<5>/Q	I0<2>/I1<5>/Q#2	   56.4103	$poly_conn
Rl137	I0<2>/I1<5>/Q#2	I0<2>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl138	WL#90	WL#91	   59.7064	$poly_conn
Rl139	WL#91	WL#92	   59.7064	$poly_conn
Rl140	I0<2>/I1<7>/Q	I0<2>/I1<7>/Q#2	   90.3330	$poly_conn
Rl141	I0<2>/I1<7>/Q#2	I0<2>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl142	I0<2>/I1<7>/QB	I0<2>/I1<7>/QB#2	   56.4103	$poly_conn
Rl143	I0<2>/I1<7>/QB#2	I0<2>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl144	WL#94	WL#95	   59.7064	$poly_conn
Rl145	WL#95	WL#96	   59.7064	$poly_conn
Rl146	I0<3>/I1<0>/QB	I0<3>/I1<0>/QB#2	   56.4103	$poly_conn
Rl147	I0<3>/I1<0>/QB	I0<3>/I1<0>/QB#3	   90.3330	$poly_conn
Rl148	I0<3>/I1<0>/Q	I0<3>/I1<0>/Q#2	   56.4103	$poly_conn
Rl149	I0<3>/I1<0>/Q#2	I0<3>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl150	WL#98	WL#99	   59.7064	$poly_conn
Rl151	WL#99	WL#100	   59.7064	$poly_conn
Rl152	I0<3>/I1<2>/Q	I0<3>/I1<2>/Q#2	   90.3330	$poly_conn
Rl153	I0<3>/I1<2>/Q#2	I0<3>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl154	I0<3>/I1<2>/QB	I0<3>/I1<2>/QB#2	   56.4103	$poly_conn
Rl155	I0<3>/I1<2>/QB#2	I0<3>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl156	WL#102	WL#103	   59.7064	$poly_conn
Rl157	WL#103	WL#104	   59.7064	$poly_conn
Rl158	I0<3>/I1<1>/QB	I0<3>/I1<1>/QB#2	   56.4103	$poly_conn
Rl159	I0<3>/I1<1>/QB	I0<3>/I1<1>/QB#3	   90.3330	$poly_conn
Rl160	I0<3>/I1<1>/Q	I0<3>/I1<1>/Q#2	   56.4103	$poly_conn
Rl161	I0<3>/I1<1>/Q#2	I0<3>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl162	WL#106	WL#107	   59.7064	$poly_conn
Rl163	WL#107	WL#108	   59.7064	$poly_conn
Rl164	I0<3>/I1<4>/Q	I0<3>/I1<4>/Q#2	   90.3330	$poly_conn
Rl165	I0<3>/I1<4>/Q#2	I0<3>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl166	I0<3>/I1<4>/QB	I0<3>/I1<4>/QB#2	   56.4103	$poly_conn
Rl167	I0<3>/I1<4>/QB#2	I0<3>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl168	WL#110	WL#111	   59.7064	$poly_conn
Rl169	WL#111	WL#112	   59.7064	$poly_conn
Rl170	I0<3>/I1<3>/QB	I0<3>/I1<3>/QB#2	   56.4103	$poly_conn
Rl171	I0<3>/I1<3>/QB	I0<3>/I1<3>/QB#3	   90.3330	$poly_conn
Rl172	I0<3>/I1<3>/Q	I0<3>/I1<3>/Q#2	   56.4103	$poly_conn
Rl173	I0<3>/I1<3>/Q#2	I0<3>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl174	WL#114	WL#115	   59.7064	$poly_conn
Rl175	WL#115	WL#116	   59.7064	$poly_conn
Rl176	I0<3>/I1<6>/Q	I0<3>/I1<6>/Q#2	   90.3330	$poly_conn
Rl177	I0<3>/I1<6>/Q#2	I0<3>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl178	I0<3>/I1<6>/QB	I0<3>/I1<6>/QB#2	   56.4103	$poly_conn
Rl179	I0<3>/I1<6>/QB#2	I0<3>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl180	WL#118	WL#119	   59.7064	$poly_conn
Rl181	WL#119	WL#120	   59.7064	$poly_conn
Rl182	I0<3>/I1<5>/QB	I0<3>/I1<5>/QB#2	   56.4103	$poly_conn
Rl183	I0<3>/I1<5>/QB	I0<3>/I1<5>/QB#3	   90.3330	$poly_conn
Rl184	I0<3>/I1<5>/Q	I0<3>/I1<5>/Q#2	   56.4103	$poly_conn
Rl185	I0<3>/I1<5>/Q#2	I0<3>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl186	WL#122	WL#123	   59.7064	$poly_conn
Rl187	WL#123	WL#124	   59.7064	$poly_conn
Rl188	I0<3>/I1<7>/Q	I0<3>/I1<7>/Q#2	   90.3330	$poly_conn
Rl189	I0<3>/I1<7>/Q#2	I0<3>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl190	I0<3>/I1<7>/QB	I0<3>/I1<7>/QB#2	   56.4103	$poly_conn
Rl191	I0<3>/I1<7>/QB#2	I0<3>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl192	WL#126	WL#127	   59.7064	$poly_conn
Rl193	WL#127	WL#128	   59.7064	$poly_conn
Rl194	I0<4>/I1<0>/QB	I0<4>/I1<0>/QB#2	   56.4103	$poly_conn
Rl195	I0<4>/I1<0>/QB	I0<4>/I1<0>/QB#3	   90.3330	$poly_conn
Rl196	I0<4>/I1<0>/Q	I0<4>/I1<0>/Q#2	   56.4103	$poly_conn
Rl197	I0<4>/I1<0>/Q#2	I0<4>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl198	WL#130	WL#131	   59.7064	$poly_conn
Rl199	WL#131	WL#132	   59.7064	$poly_conn
Rl200	I0<4>/I1<2>/Q	I0<4>/I1<2>/Q#2	   90.3330	$poly_conn
Rl201	I0<4>/I1<2>/Q#2	I0<4>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl202	I0<4>/I1<2>/QB	I0<4>/I1<2>/QB#2	   56.4103	$poly_conn
Rl203	I0<4>/I1<2>/QB#2	I0<4>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl204	WL#134	WL#135	   59.7064	$poly_conn
Rl205	WL#135	WL#136	   59.7064	$poly_conn
Rl206	I0<4>/I1<1>/QB	I0<4>/I1<1>/QB#2	   56.4103	$poly_conn
Rl207	I0<4>/I1<1>/QB	I0<4>/I1<1>/QB#3	   90.3330	$poly_conn
Rl208	I0<4>/I1<1>/Q	I0<4>/I1<1>/Q#2	   56.4103	$poly_conn
Rl209	I0<4>/I1<1>/Q#2	I0<4>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl210	WL#138	WL#139	   59.7064	$poly_conn
Rl211	WL#139	WL#140	   59.7064	$poly_conn
Rl212	I0<4>/I1<4>/Q	I0<4>/I1<4>/Q#2	   90.3330	$poly_conn
Rl213	I0<4>/I1<4>/Q#2	I0<4>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl214	I0<4>/I1<4>/QB	I0<4>/I1<4>/QB#2	   56.4103	$poly_conn
Rl215	I0<4>/I1<4>/QB#2	I0<4>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl216	WL#142	WL#143	   59.7064	$poly_conn
Rl217	WL#143	WL#144	   59.7064	$poly_conn
Rl218	I0<4>/I1<3>/QB	I0<4>/I1<3>/QB#2	   56.4103	$poly_conn
Rl219	I0<4>/I1<3>/QB	I0<4>/I1<3>/QB#3	   90.3330	$poly_conn
Rl220	I0<4>/I1<3>/Q	I0<4>/I1<3>/Q#2	   56.4103	$poly_conn
Rl221	I0<4>/I1<3>/Q#2	I0<4>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl222	WL#146	WL#147	   59.7064	$poly_conn
Rl223	WL#147	WL#148	   59.7064	$poly_conn
Rl224	I0<4>/I1<6>/Q	I0<4>/I1<6>/Q#2	   90.3330	$poly_conn
Rl225	I0<4>/I1<6>/Q#2	I0<4>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl226	I0<4>/I1<6>/QB	I0<4>/I1<6>/QB#2	   56.4103	$poly_conn
Rl227	I0<4>/I1<6>/QB#2	I0<4>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl228	WL#150	WL#151	   59.7064	$poly_conn
Rl229	WL#151	WL#152	   59.7064	$poly_conn
Rl230	I0<4>/I1<5>/QB	I0<4>/I1<5>/QB#2	   56.4103	$poly_conn
Rl231	I0<4>/I1<5>/QB	I0<4>/I1<5>/QB#3	   90.3330	$poly_conn
Rl232	I0<4>/I1<5>/Q	I0<4>/I1<5>/Q#2	   56.4103	$poly_conn
Rl233	I0<4>/I1<5>/Q#2	I0<4>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl234	WL#154	WL#155	   59.7064	$poly_conn
Rl235	WL#155	WL#156	   59.7064	$poly_conn
Rl236	I0<4>/I1<7>/Q	I0<4>/I1<7>/Q#2	   90.3330	$poly_conn
Rl237	I0<4>/I1<7>/Q#2	I0<4>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl238	I0<4>/I1<7>/QB	I0<4>/I1<7>/QB#2	   56.4103	$poly_conn
Rl239	I0<4>/I1<7>/QB#2	I0<4>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl240	WL#158	WL#159	   59.7064	$poly_conn
Rl241	WL#159	WL#160	   59.7064	$poly_conn
Rl242	I0<5>/I1<0>/QB	I0<5>/I1<0>/QB#2	   56.4103	$poly_conn
Rl243	I0<5>/I1<0>/QB	I0<5>/I1<0>/QB#3	   90.3330	$poly_conn
Rl244	I0<5>/I1<0>/Q	I0<5>/I1<0>/Q#2	   56.4103	$poly_conn
Rl245	I0<5>/I1<0>/Q#2	I0<5>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl246	WL#162	WL#163	   59.7064	$poly_conn
Rl247	WL#163	WL#164	   59.7064	$poly_conn
Rl248	I0<5>/I1<2>/Q	I0<5>/I1<2>/Q#2	   90.3330	$poly_conn
Rl249	I0<5>/I1<2>/Q#2	I0<5>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl250	I0<5>/I1<2>/QB	I0<5>/I1<2>/QB#2	   56.4103	$poly_conn
Rl251	I0<5>/I1<2>/QB#2	I0<5>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl252	WL#166	WL#167	   59.7064	$poly_conn
Rl253	WL#167	WL#168	   59.7064	$poly_conn
Rl254	I0<5>/I1<1>/QB	I0<5>/I1<1>/QB#2	   56.4103	$poly_conn
Rl255	I0<5>/I1<1>/QB	I0<5>/I1<1>/QB#3	   90.3330	$poly_conn
Rl256	I0<5>/I1<1>/Q	I0<5>/I1<1>/Q#2	   56.4103	$poly_conn
Rl257	I0<5>/I1<1>/Q#2	I0<5>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl258	WL#170	WL#171	   59.7064	$poly_conn
Rl259	WL#171	WL#172	   59.7064	$poly_conn
Rl260	I0<5>/I1<4>/Q	I0<5>/I1<4>/Q#2	   90.3330	$poly_conn
Rl261	I0<5>/I1<4>/Q#2	I0<5>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl262	I0<5>/I1<4>/QB	I0<5>/I1<4>/QB#2	   56.4103	$poly_conn
Rl263	I0<5>/I1<4>/QB#2	I0<5>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl264	WL#174	WL#175	   59.7064	$poly_conn
Rl265	WL#175	WL#176	   59.7064	$poly_conn
Rl266	I0<5>/I1<3>/QB	I0<5>/I1<3>/QB#2	   56.4103	$poly_conn
Rl267	I0<5>/I1<3>/QB	I0<5>/I1<3>/QB#3	   90.3330	$poly_conn
Rl268	I0<5>/I1<3>/Q	I0<5>/I1<3>/Q#2	   56.4103	$poly_conn
Rl269	I0<5>/I1<3>/Q#2	I0<5>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl270	WL#178	WL#179	   59.7064	$poly_conn
Rl271	WL#179	WL#180	   59.7064	$poly_conn
Rl272	I0<5>/I1<6>/Q	I0<5>/I1<6>/Q#2	   90.3330	$poly_conn
Rl273	I0<5>/I1<6>/Q#2	I0<5>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl274	I0<5>/I1<6>/QB	I0<5>/I1<6>/QB#2	   56.4103	$poly_conn
Rl275	I0<5>/I1<6>/QB#2	I0<5>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl276	WL#182	WL#183	   59.7064	$poly_conn
Rl277	WL#183	WL#184	   59.7064	$poly_conn
Rl278	I0<5>/I1<5>/QB	I0<5>/I1<5>/QB#2	   56.4103	$poly_conn
Rl279	I0<5>/I1<5>/QB	I0<5>/I1<5>/QB#3	   90.3330	$poly_conn
Rl280	I0<5>/I1<5>/Q	I0<5>/I1<5>/Q#2	   56.4103	$poly_conn
Rl281	I0<5>/I1<5>/Q#2	I0<5>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl282	WL#186	WL#187	   59.7064	$poly_conn
Rl283	WL#187	WL#188	   59.7064	$poly_conn
Rl284	I0<5>/I1<7>/Q	I0<5>/I1<7>/Q#2	   90.3330	$poly_conn
Rl285	I0<5>/I1<7>/Q#2	I0<5>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl286	I0<5>/I1<7>/QB	I0<5>/I1<7>/QB#2	   56.4103	$poly_conn
Rl287	I0<5>/I1<7>/QB#2	I0<5>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl288	WL#190	WL#191	   59.7064	$poly_conn
Rl289	WL#191	WL#192	   59.7064	$poly_conn
Rl290	I0<6>/I1<0>/QB	I0<6>/I1<0>/QB#2	   56.4103	$poly_conn
Rl291	I0<6>/I1<0>/QB	I0<6>/I1<0>/QB#3	   90.3330	$poly_conn
Rl292	I0<6>/I1<0>/Q	I0<6>/I1<0>/Q#2	   56.4103	$poly_conn
Rl293	I0<6>/I1<0>/Q#2	I0<6>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl294	WL#194	WL#195	   59.7064	$poly_conn
Rl295	WL#195	WL#196	   59.7064	$poly_conn
Rl296	I0<6>/I1<2>/Q	I0<6>/I1<2>/Q#2	   90.3330	$poly_conn
Rl297	I0<6>/I1<2>/Q#2	I0<6>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl298	I0<6>/I1<2>/QB	I0<6>/I1<2>/QB#2	   56.4103	$poly_conn
Rl299	I0<6>/I1<2>/QB#2	I0<6>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl300	WL#198	WL#199	   59.7064	$poly_conn
Rl301	WL#199	WL#200	   59.7064	$poly_conn
Rl302	I0<6>/I1<1>/QB	I0<6>/I1<1>/QB#2	   56.4103	$poly_conn
Rl303	I0<6>/I1<1>/QB	I0<6>/I1<1>/QB#3	   90.3330	$poly_conn
Rl304	I0<6>/I1<1>/Q	I0<6>/I1<1>/Q#2	   56.4103	$poly_conn
Rl305	I0<6>/I1<1>/Q#2	I0<6>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl306	WL#202	WL#203	   59.7064	$poly_conn
Rl307	WL#203	WL#204	   59.7064	$poly_conn
Rl308	I0<6>/I1<4>/Q	I0<6>/I1<4>/Q#2	   90.3330	$poly_conn
Rl309	I0<6>/I1<4>/Q#2	I0<6>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl310	I0<6>/I1<4>/QB	I0<6>/I1<4>/QB#2	   56.4103	$poly_conn
Rl311	I0<6>/I1<4>/QB#2	I0<6>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl312	WL#206	WL#207	   59.7064	$poly_conn
Rl313	WL#207	WL#208	   59.7064	$poly_conn
Rl314	I0<6>/I1<3>/QB	I0<6>/I1<3>/QB#2	   56.4103	$poly_conn
Rl315	I0<6>/I1<3>/QB	I0<6>/I1<3>/QB#3	   90.3330	$poly_conn
Rl316	I0<6>/I1<3>/Q	I0<6>/I1<3>/Q#2	   56.4103	$poly_conn
Rl317	I0<6>/I1<3>/Q#2	I0<6>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl318	WL#210	WL#211	   59.7064	$poly_conn
Rl319	WL#211	WL#212	   59.7064	$poly_conn
Rl320	I0<6>/I1<6>/Q	I0<6>/I1<6>/Q#2	   90.3330	$poly_conn
Rl321	I0<6>/I1<6>/Q#2	I0<6>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl322	I0<6>/I1<6>/QB	I0<6>/I1<6>/QB#2	   56.4103	$poly_conn
Rl323	I0<6>/I1<6>/QB#2	I0<6>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl324	WL#214	WL#215	   59.7064	$poly_conn
Rl325	WL#215	WL#216	   59.7064	$poly_conn
Rl326	I0<6>/I1<5>/QB	I0<6>/I1<5>/QB#2	   56.4103	$poly_conn
Rl327	I0<6>/I1<5>/QB	I0<6>/I1<5>/QB#3	   90.3330	$poly_conn
Rl328	I0<6>/I1<5>/Q	I0<6>/I1<5>/Q#2	   56.4103	$poly_conn
Rl329	I0<6>/I1<5>/Q#2	I0<6>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl330	WL#218	WL#219	   59.7064	$poly_conn
Rl331	WL#219	WL#220	   59.7064	$poly_conn
Rl332	I0<6>/I1<7>/Q	I0<6>/I1<7>/Q#2	   90.3330	$poly_conn
Rl333	I0<6>/I1<7>/Q#2	I0<6>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl334	I0<6>/I1<7>/QB	I0<6>/I1<7>/QB#2	   56.4103	$poly_conn
Rl335	I0<6>/I1<7>/QB#2	I0<6>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl336	WL#222	WL#223	   59.7064	$poly_conn
Rl337	WL#223	WL#224	   59.7064	$poly_conn
Rl338	I0<7>/I1<0>/QB	I0<7>/I1<0>/QB#2	   56.4103	$poly_conn
Rl339	I0<7>/I1<0>/QB	I0<7>/I1<0>/QB#3	   90.3330	$poly_conn
Rl340	I0<7>/I1<0>/Q	I0<7>/I1<0>/Q#2	   56.4103	$poly_conn
Rl341	I0<7>/I1<0>/Q#2	I0<7>/I1<0>/Q#3	   90.3330
+ $poly_conn
Rl342	WL#226	WL#227	   59.7064	$poly_conn
Rl343	WL#227	WL#228	   59.7064	$poly_conn
Rl344	I0<7>/I1<2>/Q	I0<7>/I1<2>/Q#2	   90.3330	$poly_conn
Rl345	I0<7>/I1<2>/Q#2	I0<7>/I1<2>/Q#3	   56.4103
+ $poly_conn
Rl346	I0<7>/I1<2>/QB	I0<7>/I1<2>/QB#2	   56.4103	$poly_conn
Rl347	I0<7>/I1<2>/QB#2	I0<7>/I1<2>/QB#3	   90.3330
+ $poly_conn
Rl348	WL#230	WL#231	   59.7064	$poly_conn
Rl349	WL#231	WL#232	   59.7064	$poly_conn
Rl350	I0<7>/I1<1>/QB	I0<7>/I1<1>/QB#2	   56.4103	$poly_conn
Rl351	I0<7>/I1<1>/QB	I0<7>/I1<1>/QB#3	   90.3330	$poly_conn
Rl352	I0<7>/I1<1>/Q	I0<7>/I1<1>/Q#2	   56.4103	$poly_conn
Rl353	I0<7>/I1<1>/Q#2	I0<7>/I1<1>/Q#3	   90.3330
+ $poly_conn
Rl354	WL#234	WL#235	   59.7064	$poly_conn
Rl355	WL#235	WL#236	   59.7064	$poly_conn
Rl356	I0<7>/I1<4>/Q	I0<7>/I1<4>/Q#2	   90.3330	$poly_conn
Rl357	I0<7>/I1<4>/Q#2	I0<7>/I1<4>/Q#3	   56.4103
+ $poly_conn
Rl358	I0<7>/I1<4>/QB	I0<7>/I1<4>/QB#2	   56.4103	$poly_conn
Rl359	I0<7>/I1<4>/QB#2	I0<7>/I1<4>/QB#3	   90.3330
+ $poly_conn
Rl360	WL#238	WL#239	   59.7064	$poly_conn
Rl361	WL#239	WL#240	   59.7064	$poly_conn
Rl362	I0<7>/I1<3>/QB	I0<7>/I1<3>/QB#2	   56.4103	$poly_conn
Rl363	I0<7>/I1<3>/QB	I0<7>/I1<3>/QB#3	   90.3330	$poly_conn
Rl364	I0<7>/I1<3>/Q	I0<7>/I1<3>/Q#2	   56.4103	$poly_conn
Rl365	I0<7>/I1<3>/Q#2	I0<7>/I1<3>/Q#3	   90.3330
+ $poly_conn
Rl366	WL#242	WL#243	   59.7064	$poly_conn
Rl367	WL#243	WL#244	   59.7064	$poly_conn
Rl368	I0<7>/I1<6>/Q	I0<7>/I1<6>/Q#2	   90.3330	$poly_conn
Rl369	I0<7>/I1<6>/Q#2	I0<7>/I1<6>/Q#3	   56.4103
+ $poly_conn
Rl370	I0<7>/I1<6>/QB	I0<7>/I1<6>/QB#2	   56.4103	$poly_conn
Rl371	I0<7>/I1<6>/QB#2	I0<7>/I1<6>/QB#3	   90.3330
+ $poly_conn
Rl372	WL#246	WL#247	   59.7064	$poly_conn
Rl373	WL#247	WL#248	   59.7064	$poly_conn
Rl374	I0<7>/I1<5>/QB	I0<7>/I1<5>/QB#2	   56.4103	$poly_conn
Rl375	I0<7>/I1<5>/QB	I0<7>/I1<5>/QB#3	   90.3330	$poly_conn
Rl376	I0<7>/I1<5>/Q	I0<7>/I1<5>/Q#2	   56.4103	$poly_conn
Rl377	I0<7>/I1<5>/Q#2	I0<7>/I1<5>/Q#3	   90.3330
+ $poly_conn
Rl378	WL#250	WL#251	   59.7064	$poly_conn
Rl379	WL#251	WL#252	   59.7064	$poly_conn
Rl380	I0<7>/I1<7>/Q	I0<7>/I1<7>/Q#2	   90.3330	$poly_conn
Rl381	I0<7>/I1<7>/Q#2	I0<7>/I1<7>/Q#3	   56.4103
+ $poly_conn
Rl382	I0<7>/I1<7>/QB	I0<7>/I1<7>/QB#2	   56.4103	$poly_conn
Rl383	I0<7>/I1<7>/QB#2	I0<7>/I1<7>/QB#3	   90.3330
+ $poly_conn
Rl384	WL#254	WL#255	  104.7064	$poly_conn
Rk1	WL#2	WL#9	    6.6000	$metal1_conn
Rk2	VSS#4	VSS#3	   27.3715	$metal1_conn
Rk3	VSS#6	VSS#2	   75.1654	$metal1_conn
Rk4	BL<0>#1	BL<0>#2	   81.6000	$metal1_conn
Rk5	I0<0>/I1<0>/Q#3	I0<0>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk6	I0<0>/I1<0>/Q#5	I0<0>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk7	I0<0>/I1<0>/Q#4	I0<0>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk8	VDD#1	VDD#2	   68.7306	$metal1_conn
Rk9	VDD#3	VDD#4	   31.6000	$metal1_conn
Rk10	VDD#5	VDD#6	   68.7306	$metal1_conn
Rk11	BLB<0>#3	BLB<0>#1	   75.0000	$metal1_conn
Rk12	I0<0>/I1<0>/QB#4	I0<0>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk13	I0<0>/I1<0>/QB#6	I0<0>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk14	I0<0>/I1<0>/QB#5	I0<0>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk15	WL#4	WL#13	   51.6000	$metal1_conn
Rk16	VSS#7	VSS#4	   19.0550	$metal1_conn
Rk17	VSS#11	VSS#8	   75.1654	$metal1_conn
Rk18	VSS#8	VSS#12	   75.1654	$metal1_conn
Rk19	BLB<1>#1	BLB<1>#2	   81.6000	$metal1_conn
Rk20	I0<0>/I1<2>/QB#3	I0<0>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk21	I0<0>/I1<2>/QB#5	I0<0>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk22	I0<0>/I1<2>/QB#4	I0<0>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk23	VDD#10	VDD#11	   68.7306	$metal1_conn
Rk24	VDD#12	VDD#13	   31.6000	$metal1_conn
Rk25	VDD#14	VDD#15	   68.7306	$metal1_conn
Rk26	BL<1>#1	BL<1>#2	   81.6000	$metal1_conn
Rk27	I0<0>/I1<2>/Q#4	I0<0>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk28	I0<0>/I1<2>/Q#6	I0<0>/I1<2>/Q	    0.1668	$metal1_conn
Rk29	I0<0>/I1<2>/Q#5	I0<0>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk30	WL#7	WL#17	   51.6000	$metal1_conn
Rk31	VSS#15	VSS#4	   19.0550	$metal1_conn
Rk32	VSS#17	VSS#14	   75.1654	$metal1_conn
Rk33	VSS#14	VSS#18	   75.1654	$metal1_conn
Rk34	BL<2>#1	BL<2>#2	   81.6000	$metal1_conn
Rk35	I0<0>/I1<1>/Q#3	I0<0>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk36	I0<0>/I1<1>/Q#5	I0<0>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk37	I0<0>/I1<1>/Q#4	I0<0>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk38	VDD#19	VDD#20	   68.7306	$metal1_conn
Rk39	VDD#21	VDD#22	   31.6000	$metal1_conn
Rk40	VDD#23	VDD#24	   68.7306	$metal1_conn
Rk41	BLB<2>#3	BLB<2>#1	   75.0000	$metal1_conn
Rk42	I0<0>/I1<1>/QB#4	I0<0>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk43	I0<0>/I1<1>/QB#6	I0<0>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk44	I0<0>/I1<1>/QB#5	I0<0>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk45	WL#11	WL#21	   51.6000	$metal1_conn
Rk46	VSS#19	VSS#4	   19.0550	$metal1_conn
Rk47	VSS#23	VSS#20	   75.1654	$metal1_conn
Rk48	VSS#20	VSS#24	   75.1654	$metal1_conn
Rk49	BLB<3>#1	BLB<3>#2	   81.6000	$metal1_conn
Rk50	I0<0>/I1<4>/QB#3	I0<0>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk51	I0<0>/I1<4>/QB#5	I0<0>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk52	I0<0>/I1<4>/QB#4	I0<0>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk53	VDD#28	VDD#29	   68.7306	$metal1_conn
Rk54	VDD#30	VDD#31	   31.6000	$metal1_conn
Rk55	VDD#32	VDD#33	   68.7306	$metal1_conn
Rk56	BL<3>#1	BL<3>#2	   81.6000	$metal1_conn
Rk57	I0<0>/I1<4>/Q#4	I0<0>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk58	I0<0>/I1<4>/Q#6	I0<0>/I1<4>/Q	    0.1668	$metal1_conn
Rk59	I0<0>/I1<4>/Q#5	I0<0>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk60	WL#15	WL#25	   51.6000	$metal1_conn
Rk61	VSS#27	VSS#4	   19.0550	$metal1_conn
Rk62	VSS#29	VSS#26	   75.1654	$metal1_conn
Rk63	VSS#26	VSS#30	   75.1654	$metal1_conn
Rk64	BL<4>#1	BL<4>#2	   81.6000	$metal1_conn
Rk65	I0<0>/I1<3>/Q#3	I0<0>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk66	I0<0>/I1<3>/Q#5	I0<0>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk67	I0<0>/I1<3>/Q#4	I0<0>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk68	VDD#37	VDD#38	   68.7306	$metal1_conn
Rk69	VDD#39	VDD#40	   31.6000	$metal1_conn
Rk70	VDD#41	VDD#42	   68.7306	$metal1_conn
Rk71	BLB<4>#3	BLB<4>#1	   75.0000	$metal1_conn
Rk72	I0<0>/I1<3>/QB#4	I0<0>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk73	I0<0>/I1<3>/QB#6	I0<0>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk74	I0<0>/I1<3>/QB#5	I0<0>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk75	WL#19	WL#29	   51.6000	$metal1_conn
Rk76	VSS#31	VSS#4	   19.0550	$metal1_conn
Rk77	VSS#35	VSS#32	   75.1654	$metal1_conn
Rk78	VSS#32	VSS#36	   75.1654	$metal1_conn
Rk79	BLB<5>#1	BLB<5>#2	   81.6000	$metal1_conn
Rk80	I0<0>/I1<6>/QB#3	I0<0>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk81	I0<0>/I1<6>/QB#5	I0<0>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk82	I0<0>/I1<6>/QB#4	I0<0>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk83	VDD#46	VDD#47	   68.7306	$metal1_conn
Rk84	VDD#48	VDD#49	   31.6000	$metal1_conn
Rk85	VDD#50	VDD#51	   68.7306	$metal1_conn
Rk86	BL<5>#1	BL<5>#2	   81.6000	$metal1_conn
Rk87	I0<0>/I1<6>/Q#4	I0<0>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk88	I0<0>/I1<6>/Q#6	I0<0>/I1<6>/Q	    0.1668	$metal1_conn
Rk89	I0<0>/I1<6>/Q#5	I0<0>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk90	WL#23	WL#33	   51.6000	$metal1_conn
Rk91	VSS#39	VSS#4	   19.0550	$metal1_conn
Rk92	VSS#41	VSS#38	   75.1654	$metal1_conn
Rk93	VSS#38	VSS#42	   75.1654	$metal1_conn
Rk94	BL<6>#1	BL<6>#2	   81.6000	$metal1_conn
Rk95	I0<0>/I1<5>/Q#3	I0<0>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk96	I0<0>/I1<5>/Q#5	I0<0>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk97	I0<0>/I1<5>/Q#4	I0<0>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk98	VDD#55	VDD#56	   68.7306	$metal1_conn
Rk99	VDD#57	VDD#58	   31.6000	$metal1_conn
Rk100	VDD#59	VDD#60	   68.7306	$metal1_conn
Rk101	BLB<6>#3	BLB<6>#1	   75.0000	$metal1_conn
Rk102	I0<0>/I1<5>/QB#4	I0<0>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk103	I0<0>/I1<5>/QB#6	I0<0>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk104	I0<0>/I1<5>/QB#5	I0<0>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk105	WL#27	WL#37	   51.6000	$metal1_conn
Rk106	VSS#43	VSS#4	   19.0550	$metal1_conn
Rk107	VSS#47	VSS#44	   75.1654	$metal1_conn
Rk108	VSS#44	VSS#48	   75.1654	$metal1_conn
Rk109	BLB<7>#1	BLB<7>#2	   81.6000	$metal1_conn
Rk110	I0<0>/I1<7>/QB#3	I0<0>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk111	I0<0>/I1<7>/QB#5	I0<0>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk112	I0<0>/I1<7>/QB#4	I0<0>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk113	VDD#64	VDD#65	   68.7306	$metal1_conn
Rk114	VDD#66	VDD#67	   31.6000	$metal1_conn
Rk115	VDD#68	VDD#69	   68.7306	$metal1_conn
Rk116	BL<7>#1	BL<7>#2	   81.6000	$metal1_conn
Rk117	I0<0>/I1<7>/Q#4	I0<0>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk118	I0<0>/I1<7>/Q#6	I0<0>/I1<7>/Q	    0.1668	$metal1_conn
Rk119	I0<0>/I1<7>/Q#5	I0<0>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk120	WL#31	WL#41	   51.6000	$metal1_conn
Rk121	VSS#51	VSS#4	   19.0550	$metal1_conn
Rk122	VSS#53	VSS#50	   75.1654	$metal1_conn
Rk123	VSS#50	VSS#54	   75.1654	$metal1_conn
Rk124	BL<8>#1	BL<8>#2	   81.6000	$metal1_conn
Rk125	I0<1>/I1<0>/Q#3	I0<1>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk126	I0<1>/I1<0>/Q#5	I0<1>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk127	I0<1>/I1<0>/Q#4	I0<1>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk128	VDD#73	VDD#74	   68.7306	$metal1_conn
Rk129	VDD#75	VDD#76	   31.6000	$metal1_conn
Rk130	VDD#77	VDD#78	   68.7306	$metal1_conn
Rk131	BLB<8>#3	BLB<8>#1	   75.0000	$metal1_conn
Rk132	I0<1>/I1<0>/QB#4	I0<1>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk133	I0<1>/I1<0>/QB#6	I0<1>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk134	I0<1>/I1<0>/QB#5	I0<1>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk135	WL#35	WL#45	   51.6000	$metal1_conn
Rk136	VSS#55	VSS#4	   19.0550	$metal1_conn
Rk137	VSS#59	VSS#56	   75.1654	$metal1_conn
Rk138	VSS#56	VSS#60	   75.1654	$metal1_conn
Rk139	BLB<9>#1	BLB<9>#2	   81.6000	$metal1_conn
Rk140	I0<1>/I1<2>/QB#3	I0<1>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk141	I0<1>/I1<2>/QB#5	I0<1>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk142	I0<1>/I1<2>/QB#4	I0<1>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk143	VDD#82	VDD#83	   68.7306	$metal1_conn
Rk144	VDD#84	VDD#85	   31.6000	$metal1_conn
Rk145	VDD#86	VDD#87	   68.7306	$metal1_conn
Rk146	BL<9>#1	BL<9>#2	   81.6000	$metal1_conn
Rk147	I0<1>/I1<2>/Q#4	I0<1>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk148	I0<1>/I1<2>/Q#6	I0<1>/I1<2>/Q	    0.1668	$metal1_conn
Rk149	I0<1>/I1<2>/Q#5	I0<1>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk150	WL#39	WL#49	   51.6000	$metal1_conn
Rk151	VSS#63	VSS#4	   19.0550	$metal1_conn
Rk152	VSS#65	VSS#62	   75.1654	$metal1_conn
Rk153	VSS#62	VSS#66	   75.1654	$metal1_conn
Rk154	BL<10>#1	BL<10>#2	   81.6000	$metal1_conn
Rk155	I0<1>/I1<1>/Q#3	I0<1>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk156	I0<1>/I1<1>/Q#5	I0<1>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk157	I0<1>/I1<1>/Q#4	I0<1>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk158	VDD#91	VDD#92	   68.7306	$metal1_conn
Rk159	VDD#93	VDD#94	   31.6000	$metal1_conn
Rk160	VDD#95	VDD#96	   68.7306	$metal1_conn
Rk161	BLB<10>#3	BLB<10>#1	   75.0000	$metal1_conn
Rk162	I0<1>/I1<1>/QB#4	I0<1>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk163	I0<1>/I1<1>/QB#6	I0<1>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk164	I0<1>/I1<1>/QB#5	I0<1>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk165	WL#43	WL#53	   51.6000	$metal1_conn
Rk166	VSS#67	VSS#4	   19.0550	$metal1_conn
Rk167	VSS#71	VSS#68	   75.1654	$metal1_conn
Rk168	VSS#68	VSS#72	   75.1654	$metal1_conn
Rk169	BLB<11>#1	BLB<11>#2	   81.6000	$metal1_conn
Rk170	I0<1>/I1<4>/QB#3	I0<1>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk171	I0<1>/I1<4>/QB#5	I0<1>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk172	I0<1>/I1<4>/QB#4	I0<1>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk173	VDD#100	VDD#101	   68.7306	$metal1_conn
Rk174	VDD#102	VDD#103	   31.6000	$metal1_conn
Rk175	VDD#104	VDD#105	   68.7306	$metal1_conn
Rk176	BL<11>#1	BL<11>#2	   81.6000	$metal1_conn
Rk177	I0<1>/I1<4>/Q#4	I0<1>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk178	I0<1>/I1<4>/Q#6	I0<1>/I1<4>/Q	    0.1668	$metal1_conn
Rk179	I0<1>/I1<4>/Q#5	I0<1>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk180	WL#47	WL#57	   51.6000	$metal1_conn
Rk181	VSS#75	VSS#4	   19.0550	$metal1_conn
Rk182	VSS#77	VSS#74	   75.1654	$metal1_conn
Rk183	VSS#74	VSS#78	   75.1654	$metal1_conn
Rk184	BL<12>#1	BL<12>#2	   81.6000	$metal1_conn
Rk185	I0<1>/I1<3>/Q#3	I0<1>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk186	I0<1>/I1<3>/Q#5	I0<1>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk187	I0<1>/I1<3>/Q#4	I0<1>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk188	VDD#109	VDD#110	   68.7306	$metal1_conn
Rk189	VDD#111	VDD#112	   31.6000	$metal1_conn
Rk190	VDD#113	VDD#114	   68.7306	$metal1_conn
Rk191	BLB<12>#3	BLB<12>#1	   75.0000	$metal1_conn
Rk192	I0<1>/I1<3>/QB#4	I0<1>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk193	I0<1>/I1<3>/QB#6	I0<1>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk194	I0<1>/I1<3>/QB#5	I0<1>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk195	WL#51	WL#61	   51.6000	$metal1_conn
Rk196	VSS#79	VSS#4	   19.0550	$metal1_conn
Rk197	VSS#83	VSS#80	   75.1654	$metal1_conn
Rk198	VSS#80	VSS#84	   75.1654	$metal1_conn
Rk199	BLB<13>#1	BLB<13>#2	   81.6000	$metal1_conn
Rk200	I0<1>/I1<6>/QB#3	I0<1>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk201	I0<1>/I1<6>/QB#5	I0<1>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk202	I0<1>/I1<6>/QB#4	I0<1>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk203	VDD#118	VDD#119	   68.7306	$metal1_conn
Rk204	VDD#120	VDD#121	   31.6000	$metal1_conn
Rk205	VDD#122	VDD#123	   68.7306	$metal1_conn
Rk206	BL<13>#1	BL<13>#2	   81.6000	$metal1_conn
Rk207	I0<1>/I1<6>/Q#4	I0<1>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk208	I0<1>/I1<6>/Q#6	I0<1>/I1<6>/Q	    0.1668	$metal1_conn
Rk209	I0<1>/I1<6>/Q#5	I0<1>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk210	WL#55	WL#65	   51.6000	$metal1_conn
Rk211	VSS#87	VSS#4	   19.0550	$metal1_conn
Rk212	VSS#89	VSS#86	   75.1654	$metal1_conn
Rk213	VSS#86	VSS#90	   75.1654	$metal1_conn
Rk214	BL<14>#1	BL<14>#2	   81.6000	$metal1_conn
Rk215	I0<1>/I1<5>/Q#3	I0<1>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk216	I0<1>/I1<5>/Q#5	I0<1>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk217	I0<1>/I1<5>/Q#4	I0<1>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk218	VDD#127	VDD#128	   68.7306	$metal1_conn
Rk219	VDD#129	VDD#130	   31.6000	$metal1_conn
Rk220	VDD#131	VDD#132	   68.7306	$metal1_conn
Rk221	BLB<14>#3	BLB<14>#1	   75.0000	$metal1_conn
Rk222	I0<1>/I1<5>/QB#4	I0<1>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk223	I0<1>/I1<5>/QB#6	I0<1>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk224	I0<1>/I1<5>/QB#5	I0<1>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk225	WL#59	WL#69	   51.6000	$metal1_conn
Rk226	VSS#91	VSS#4	   19.0550	$metal1_conn
Rk227	VSS#95	VSS#92	   75.1654	$metal1_conn
Rk228	VSS#92	VSS#96	   75.1654	$metal1_conn
Rk229	BLB<15>#1	BLB<15>#2	   81.6000	$metal1_conn
Rk230	I0<1>/I1<7>/QB#3	I0<1>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk231	I0<1>/I1<7>/QB#5	I0<1>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk232	I0<1>/I1<7>/QB#4	I0<1>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk233	VDD#136	VDD#137	   68.7306	$metal1_conn
Rk234	VDD#138	VDD#139	   31.6000	$metal1_conn
Rk235	VDD#140	VDD#141	   68.7306	$metal1_conn
Rk236	BL<15>#1	BL<15>#2	   81.6000	$metal1_conn
Rk237	I0<1>/I1<7>/Q#4	I0<1>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk238	I0<1>/I1<7>/Q#6	I0<1>/I1<7>/Q	    0.1668	$metal1_conn
Rk239	I0<1>/I1<7>/Q#5	I0<1>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk240	WL#63	WL#73	   51.6000	$metal1_conn
Rk241	VSS#99	VSS#4	   19.0550	$metal1_conn
Rk242	VSS#101	VSS#98	   75.1654	$metal1_conn
Rk243	VSS#98	VSS#102	   75.1654	$metal1_conn
Rk244	BL<16>#1	BL<16>#2	   81.6000	$metal1_conn
Rk245	I0<2>/I1<0>/Q#3	I0<2>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk246	I0<2>/I1<0>/Q#5	I0<2>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk247	I0<2>/I1<0>/Q#4	I0<2>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk248	VDD#145	VDD#146	   68.7306	$metal1_conn
Rk249	VDD#147	VDD#148	   31.6000	$metal1_conn
Rk250	VDD#149	VDD#150	   68.7306	$metal1_conn
Rk251	BLB<16>#3	BLB<16>#1	   75.0000	$metal1_conn
Rk252	I0<2>/I1<0>/QB#4	I0<2>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk253	I0<2>/I1<0>/QB#6	I0<2>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk254	I0<2>/I1<0>/QB#5	I0<2>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk255	WL#67	WL#77	   51.6000	$metal1_conn
Rk256	VSS#103	VSS#4	   19.0550	$metal1_conn
Rk257	VSS#107	VSS#104	   75.1654	$metal1_conn
Rk258	VSS#104	VSS#108	   75.1654	$metal1_conn
Rk259	BLB<17>#1	BLB<17>#2	   81.6000	$metal1_conn
Rk260	I0<2>/I1<2>/QB#3	I0<2>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk261	I0<2>/I1<2>/QB#5	I0<2>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk262	I0<2>/I1<2>/QB#4	I0<2>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk263	VDD#154	VDD#155	   68.7306	$metal1_conn
Rk264	VDD#156	VDD#157	   31.6000	$metal1_conn
Rk265	VDD#158	VDD#159	   68.7306	$metal1_conn
Rk266	BL<17>#1	BL<17>#2	   81.6000	$metal1_conn
Rk267	I0<2>/I1<2>/Q#4	I0<2>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk268	I0<2>/I1<2>/Q#6	I0<2>/I1<2>/Q	    0.1668	$metal1_conn
Rk269	I0<2>/I1<2>/Q#5	I0<2>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk270	WL#71	WL#81	   51.6000	$metal1_conn
Rk271	VSS#111	VSS#4	   19.0550	$metal1_conn
Rk272	VSS#113	VSS#110	   75.1654	$metal1_conn
Rk273	VSS#110	VSS#114	   75.1654	$metal1_conn
Rk274	BL<18>#1	BL<18>#2	   81.6000	$metal1_conn
Rk275	I0<2>/I1<1>/Q#3	I0<2>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk276	I0<2>/I1<1>/Q#5	I0<2>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk277	I0<2>/I1<1>/Q#4	I0<2>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk278	VDD#163	VDD#164	   68.7306	$metal1_conn
Rk279	VDD#165	VDD#166	   31.6000	$metal1_conn
Rk280	VDD#167	VDD#168	   68.7306	$metal1_conn
Rk281	BLB<18>#3	BLB<18>#1	   75.0000	$metal1_conn
Rk282	I0<2>/I1<1>/QB#4	I0<2>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk283	I0<2>/I1<1>/QB#6	I0<2>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk284	I0<2>/I1<1>/QB#5	I0<2>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk285	WL#75	WL#85	   51.6000	$metal1_conn
Rk286	VSS#115	VSS#4	   19.0550	$metal1_conn
Rk287	VSS#119	VSS#116	   75.1654	$metal1_conn
Rk288	VSS#116	VSS#120	   75.1654	$metal1_conn
Rk289	BLB<19>#1	BLB<19>#2	   81.6000	$metal1_conn
Rk290	I0<2>/I1<4>/QB#3	I0<2>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk291	I0<2>/I1<4>/QB#5	I0<2>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk292	I0<2>/I1<4>/QB#4	I0<2>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk293	VDD#172	VDD#173	   68.7306	$metal1_conn
Rk294	VDD#174	VDD#175	   31.6000	$metal1_conn
Rk295	VDD#176	VDD#177	   68.7306	$metal1_conn
Rk296	BL<19>#1	BL<19>#2	   81.6000	$metal1_conn
Rk297	I0<2>/I1<4>/Q#4	I0<2>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk298	I0<2>/I1<4>/Q#6	I0<2>/I1<4>/Q	    0.1668	$metal1_conn
Rk299	I0<2>/I1<4>/Q#5	I0<2>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk300	WL#79	WL#89	   51.6000	$metal1_conn
Rk301	VSS#123	VSS#4	   19.0550	$metal1_conn
Rk302	VSS#125	VSS#122	   75.1654	$metal1_conn
Rk303	VSS#122	VSS#126	   75.1654	$metal1_conn
Rk304	BL<20>#1	BL<20>#2	   81.6000	$metal1_conn
Rk305	I0<2>/I1<3>/Q#3	I0<2>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk306	I0<2>/I1<3>/Q#5	I0<2>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk307	I0<2>/I1<3>/Q#4	I0<2>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk308	VDD#181	VDD#182	   68.7306	$metal1_conn
Rk309	VDD#183	VDD#184	   31.6000	$metal1_conn
Rk310	VDD#185	VDD#186	   68.7306	$metal1_conn
Rk311	BLB<20>#3	BLB<20>#1	   75.0000	$metal1_conn
Rk312	I0<2>/I1<3>/QB#4	I0<2>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk313	I0<2>/I1<3>/QB#6	I0<2>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk314	I0<2>/I1<3>/QB#5	I0<2>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk315	WL#83	WL#93	   51.6000	$metal1_conn
Rk316	VSS#127	VSS#4	   19.0550	$metal1_conn
Rk317	VSS#131	VSS#128	   75.1654	$metal1_conn
Rk318	VSS#128	VSS#132	   75.1654	$metal1_conn
Rk319	BLB<21>#1	BLB<21>#2	   81.6000	$metal1_conn
Rk320	I0<2>/I1<6>/QB#3	I0<2>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk321	I0<2>/I1<6>/QB#5	I0<2>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk322	I0<2>/I1<6>/QB#4	I0<2>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk323	VDD#190	VDD#191	   68.7306	$metal1_conn
Rk324	VDD#192	VDD#193	   31.6000	$metal1_conn
Rk325	VDD#194	VDD#195	   68.7306	$metal1_conn
Rk326	BL<21>#1	BL<21>#2	   81.6000	$metal1_conn
Rk327	I0<2>/I1<6>/Q#4	I0<2>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk328	I0<2>/I1<6>/Q#6	I0<2>/I1<6>/Q	    0.1668	$metal1_conn
Rk329	I0<2>/I1<6>/Q#5	I0<2>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk330	WL#87	WL#97	   51.6000	$metal1_conn
Rk331	VSS#135	VSS#4	   19.0550	$metal1_conn
Rk332	VSS#137	VSS#134	   75.1654	$metal1_conn
Rk333	VSS#134	VSS#138	   75.1654	$metal1_conn
Rk334	BL<22>#1	BL<22>#2	   81.6000	$metal1_conn
Rk335	I0<2>/I1<5>/Q#3	I0<2>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk336	I0<2>/I1<5>/Q#5	I0<2>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk337	I0<2>/I1<5>/Q#4	I0<2>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk338	VDD#199	VDD#200	   68.7306	$metal1_conn
Rk339	VDD#201	VDD#202	   31.6000	$metal1_conn
Rk340	VDD#203	VDD#204	   68.7306	$metal1_conn
Rk341	BLB<22>#3	BLB<22>#1	   75.0000	$metal1_conn
Rk342	I0<2>/I1<5>/QB#4	I0<2>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk343	I0<2>/I1<5>/QB#6	I0<2>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk344	I0<2>/I1<5>/QB#5	I0<2>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk345	WL#91	WL#101	   51.6000	$metal1_conn
Rk346	VSS#139	VSS#4	   19.0550	$metal1_conn
Rk347	VSS#143	VSS#140	   75.1654	$metal1_conn
Rk348	VSS#140	VSS#144	   75.1654	$metal1_conn
Rk349	BLB<23>#1	BLB<23>#2	   81.6000	$metal1_conn
Rk350	I0<2>/I1<7>/QB#3	I0<2>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk351	I0<2>/I1<7>/QB#5	I0<2>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk352	I0<2>/I1<7>/QB#4	I0<2>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk353	VDD#208	VDD#209	   68.7306	$metal1_conn
Rk354	VDD#210	VDD#211	   31.6000	$metal1_conn
Rk355	VDD#212	VDD#213	   68.7306	$metal1_conn
Rk356	BL<23>#1	BL<23>#2	   81.6000	$metal1_conn
Rk357	I0<2>/I1<7>/Q#4	I0<2>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk358	I0<2>/I1<7>/Q#6	I0<2>/I1<7>/Q	    0.1668	$metal1_conn
Rk359	I0<2>/I1<7>/Q#5	I0<2>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk360	WL#95	WL#105	   51.6000	$metal1_conn
Rk361	VSS#147	VSS#4	   19.0550	$metal1_conn
Rk362	VSS#149	VSS#146	   75.1654	$metal1_conn
Rk363	VSS#146	VSS#150	   75.1654	$metal1_conn
Rk364	BL<24>#1	BL<24>#2	   81.6000	$metal1_conn
Rk365	I0<3>/I1<0>/Q#3	I0<3>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk366	I0<3>/I1<0>/Q#5	I0<3>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk367	I0<3>/I1<0>/Q#4	I0<3>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk368	VDD#217	VDD#218	   68.7306	$metal1_conn
Rk369	VDD#219	VDD#220	   31.6000	$metal1_conn
Rk370	VDD#221	VDD#222	   68.7306	$metal1_conn
Rk371	BLB<24>#3	BLB<24>#1	   75.0000	$metal1_conn
Rk372	I0<3>/I1<0>/QB#4	I0<3>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk373	I0<3>/I1<0>/QB#6	I0<3>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk374	I0<3>/I1<0>/QB#5	I0<3>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk375	WL#99	WL#109	   51.6000	$metal1_conn
Rk376	VSS#151	VSS#4	   19.0550	$metal1_conn
Rk377	VSS#155	VSS#152	   75.1654	$metal1_conn
Rk378	VSS#152	VSS#156	   75.1654	$metal1_conn
Rk379	BLB<25>#1	BLB<25>#2	   81.6000	$metal1_conn
Rk380	I0<3>/I1<2>/QB#3	I0<3>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk381	I0<3>/I1<2>/QB#5	I0<3>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk382	I0<3>/I1<2>/QB#4	I0<3>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk383	VDD#226	VDD#227	   68.7306	$metal1_conn
Rk384	VDD#228	VDD#229	   31.6000	$metal1_conn
Rk385	VDD#230	VDD#231	   68.7306	$metal1_conn
Rk386	BL<25>#1	BL<25>#2	   81.6000	$metal1_conn
Rk387	I0<3>/I1<2>/Q#4	I0<3>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk388	I0<3>/I1<2>/Q#6	I0<3>/I1<2>/Q	    0.1668	$metal1_conn
Rk389	I0<3>/I1<2>/Q#5	I0<3>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk390	WL#103	WL#113	   51.6000	$metal1_conn
Rk391	VSS#159	VSS#4	   19.0550	$metal1_conn
Rk392	VSS#161	VSS#158	   75.1654	$metal1_conn
Rk393	VSS#158	VSS#162	   75.1654	$metal1_conn
Rk394	BL<26>#1	BL<26>#2	   81.6000	$metal1_conn
Rk395	I0<3>/I1<1>/Q#3	I0<3>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk396	I0<3>/I1<1>/Q#5	I0<3>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk397	I0<3>/I1<1>/Q#4	I0<3>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk398	VDD#235	VDD#236	   68.7306	$metal1_conn
Rk399	VDD#237	VDD#238	   31.6000	$metal1_conn
Rk400	VDD#239	VDD#240	   68.7306	$metal1_conn
Rk401	BLB<26>#3	BLB<26>#1	   75.0000	$metal1_conn
Rk402	I0<3>/I1<1>/QB#4	I0<3>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk403	I0<3>/I1<1>/QB#6	I0<3>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk404	I0<3>/I1<1>/QB#5	I0<3>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk405	WL#107	WL#117	   51.6000	$metal1_conn
Rk406	VSS#163	VSS#4	   19.0550	$metal1_conn
Rk407	VSS#167	VSS#164	   75.1654	$metal1_conn
Rk408	VSS#164	VSS#168	   75.1654	$metal1_conn
Rk409	BLB<27>#1	BLB<27>#2	   81.6000	$metal1_conn
Rk410	I0<3>/I1<4>/QB#3	I0<3>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk411	I0<3>/I1<4>/QB#5	I0<3>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk412	I0<3>/I1<4>/QB#4	I0<3>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk413	VDD#244	VDD#245	   68.7306	$metal1_conn
Rk414	VDD#246	VDD#247	   31.6000	$metal1_conn
Rk415	VDD#248	VDD#249	   68.7306	$metal1_conn
Rk416	BL<27>#1	BL<27>#2	   81.6000	$metal1_conn
Rk417	I0<3>/I1<4>/Q#4	I0<3>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk418	I0<3>/I1<4>/Q#6	I0<3>/I1<4>/Q	    0.1668	$metal1_conn
Rk419	I0<3>/I1<4>/Q#5	I0<3>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk420	WL#111	WL#121	   51.6000	$metal1_conn
Rk421	VSS#171	VSS#4	   19.0550	$metal1_conn
Rk422	VSS#173	VSS#170	   75.1654	$metal1_conn
Rk423	VSS#170	VSS#174	   75.1654	$metal1_conn
Rk424	BL<28>#1	BL<28>#2	   81.6000	$metal1_conn
Rk425	I0<3>/I1<3>/Q#3	I0<3>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk426	I0<3>/I1<3>/Q#5	I0<3>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk427	I0<3>/I1<3>/Q#4	I0<3>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk428	VDD#253	VDD#254	   68.7306	$metal1_conn
Rk429	VDD#255	VDD#256	   31.6000	$metal1_conn
Rk430	VDD#257	VDD#258	   68.7306	$metal1_conn
Rk431	BLB<28>#3	BLB<28>#1	   75.0000	$metal1_conn
Rk432	I0<3>/I1<3>/QB#4	I0<3>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk433	I0<3>/I1<3>/QB#6	I0<3>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk434	I0<3>/I1<3>/QB#5	I0<3>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk435	WL#115	WL#125	   51.6000	$metal1_conn
Rk436	VSS#175	VSS#4	   19.0550	$metal1_conn
Rk437	VSS#179	VSS#176	   75.1654	$metal1_conn
Rk438	VSS#176	VSS#180	   75.1654	$metal1_conn
Rk439	BLB<29>#1	BLB<29>#2	   81.6000	$metal1_conn
Rk440	I0<3>/I1<6>/QB#3	I0<3>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk441	I0<3>/I1<6>/QB#5	I0<3>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk442	I0<3>/I1<6>/QB#4	I0<3>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk443	VDD#262	VDD#263	   68.7306	$metal1_conn
Rk444	VDD#264	VDD#265	   31.6000	$metal1_conn
Rk445	VDD#266	VDD#267	   68.7306	$metal1_conn
Rk446	BL<29>#1	BL<29>#2	   81.6000	$metal1_conn
Rk447	I0<3>/I1<6>/Q#4	I0<3>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk448	I0<3>/I1<6>/Q#6	I0<3>/I1<6>/Q	    0.1668	$metal1_conn
Rk449	I0<3>/I1<6>/Q#5	I0<3>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk450	WL#119	WL#129	   51.6000	$metal1_conn
Rk451	VSS#183	VSS#4	   19.0550	$metal1_conn
Rk452	VSS#185	VSS#182	   75.1654	$metal1_conn
Rk453	VSS#182	VSS#186	   75.1654	$metal1_conn
Rk454	BL<30>#1	BL<30>#2	   81.6000	$metal1_conn
Rk455	I0<3>/I1<5>/Q#3	I0<3>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk456	I0<3>/I1<5>/Q#5	I0<3>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk457	I0<3>/I1<5>/Q#4	I0<3>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk458	VDD#271	VDD#272	   68.7306	$metal1_conn
Rk459	VDD#273	VDD#274	   31.6000	$metal1_conn
Rk460	VDD#275	VDD#276	   68.7306	$metal1_conn
Rk461	BLB<30>#3	BLB<30>#1	   75.0000	$metal1_conn
Rk462	I0<3>/I1<5>/QB#4	I0<3>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk463	I0<3>/I1<5>/QB#6	I0<3>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk464	I0<3>/I1<5>/QB#5	I0<3>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk465	WL#123	WL#133	   51.6000	$metal1_conn
Rk466	VSS#187	VSS#4	   19.0550	$metal1_conn
Rk467	VSS#191	VSS#188	   75.1654	$metal1_conn
Rk468	VSS#188	VSS#192	   75.1654	$metal1_conn
Rk469	BLB<31>#1	BLB<31>#2	   81.6000	$metal1_conn
Rk470	I0<3>/I1<7>/QB#3	I0<3>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk471	I0<3>/I1<7>/QB#5	I0<3>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk472	I0<3>/I1<7>/QB#4	I0<3>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk473	VDD#280	VDD#281	   68.7306	$metal1_conn
Rk474	VDD#282	VDD#283	   31.6000	$metal1_conn
Rk475	VDD#284	VDD#285	   68.7306	$metal1_conn
Rk476	BL<31>#1	BL<31>#2	   81.6000	$metal1_conn
Rk477	I0<3>/I1<7>/Q#4	I0<3>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk478	I0<3>/I1<7>/Q#6	I0<3>/I1<7>/Q	    0.1668	$metal1_conn
Rk479	I0<3>/I1<7>/Q#5	I0<3>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk480	WL#127	WL#137	   51.6000	$metal1_conn
Rk481	VSS#195	VSS#4	   19.0550	$metal1_conn
Rk482	VSS#197	VSS#194	   75.1654	$metal1_conn
Rk483	VSS#194	VSS#198	   75.1654	$metal1_conn
Rk484	BL<32>#1	BL<32>#2	   81.6000	$metal1_conn
Rk485	I0<4>/I1<0>/Q#3	I0<4>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk486	I0<4>/I1<0>/Q#5	I0<4>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk487	I0<4>/I1<0>/Q#4	I0<4>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk488	VDD#289	VDD#290	   68.7306	$metal1_conn
Rk489	VDD#291	VDD#292	   31.6000	$metal1_conn
Rk490	VDD#293	VDD#294	   68.7306	$metal1_conn
Rk491	BLB<32>#3	BLB<32>#1	   75.0000	$metal1_conn
Rk492	I0<4>/I1<0>/QB#4	I0<4>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk493	I0<4>/I1<0>/QB#6	I0<4>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk494	I0<4>/I1<0>/QB#5	I0<4>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk495	WL#131	WL#141	   51.6000	$metal1_conn
Rk496	VSS#199	VSS#4	   19.0550	$metal1_conn
Rk497	VSS#203	VSS#200	   75.1654	$metal1_conn
Rk498	VSS#200	VSS#204	   75.1654	$metal1_conn
Rk499	BLB<33>#1	BLB<33>#2	   81.6000	$metal1_conn
Rk500	I0<4>/I1<2>/QB#3	I0<4>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk501	I0<4>/I1<2>/QB#5	I0<4>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk502	I0<4>/I1<2>/QB#4	I0<4>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk503	VDD#298	VDD#299	   68.7306	$metal1_conn
Rk504	VDD#300	VDD#301	   31.6000	$metal1_conn
Rk505	VDD#302	VDD#303	   68.7306	$metal1_conn
Rk506	BL<33>#1	BL<33>#2	   81.6000	$metal1_conn
Rk507	I0<4>/I1<2>/Q#4	I0<4>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk508	I0<4>/I1<2>/Q#6	I0<4>/I1<2>/Q	    0.1668	$metal1_conn
Rk509	I0<4>/I1<2>/Q#5	I0<4>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk510	WL#135	WL#145	   51.6000	$metal1_conn
Rk511	VSS#207	VSS#4	   19.0550	$metal1_conn
Rk512	VSS#209	VSS#206	   75.1654	$metal1_conn
Rk513	VSS#206	VSS#210	   75.1654	$metal1_conn
Rk514	BL<34>#1	BL<34>#2	   81.6000	$metal1_conn
Rk515	I0<4>/I1<1>/Q#3	I0<4>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk516	I0<4>/I1<1>/Q#5	I0<4>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk517	I0<4>/I1<1>/Q#4	I0<4>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk518	VDD#307	VDD#308	   68.7306	$metal1_conn
Rk519	VDD#309	VDD#310	   31.6000	$metal1_conn
Rk520	VDD#311	VDD#312	   68.7306	$metal1_conn
Rk521	BLB<34>#3	BLB<34>#1	   75.0000	$metal1_conn
Rk522	I0<4>/I1<1>/QB#4	I0<4>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk523	I0<4>/I1<1>/QB#6	I0<4>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk524	I0<4>/I1<1>/QB#5	I0<4>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk525	WL#139	WL#149	   51.6000	$metal1_conn
Rk526	VSS#211	VSS#4	   19.0550	$metal1_conn
Rk527	VSS#215	VSS#212	   75.1654	$metal1_conn
Rk528	VSS#212	VSS#216	   75.1654	$metal1_conn
Rk529	BLB<35>#1	BLB<35>#2	   81.6000	$metal1_conn
Rk530	I0<4>/I1<4>/QB#3	I0<4>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk531	I0<4>/I1<4>/QB#5	I0<4>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk532	I0<4>/I1<4>/QB#4	I0<4>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk533	VDD#316	VDD#317	   68.7306	$metal1_conn
Rk534	VDD#318	VDD#319	   31.6000	$metal1_conn
Rk535	VDD#320	VDD#321	   68.7306	$metal1_conn
Rk536	BL<35>#1	BL<35>#2	   81.6000	$metal1_conn
Rk537	I0<4>/I1<4>/Q#4	I0<4>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk538	I0<4>/I1<4>/Q#6	I0<4>/I1<4>/Q	    0.1668	$metal1_conn
Rk539	I0<4>/I1<4>/Q#5	I0<4>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk540	WL#143	WL#153	   51.6000	$metal1_conn
Rk541	VSS#219	VSS#4	   19.0550	$metal1_conn
Rk542	VSS#221	VSS#218	   75.1654	$metal1_conn
Rk543	VSS#218	VSS#222	   75.1654	$metal1_conn
Rk544	BL<36>#1	BL<36>#2	   81.6000	$metal1_conn
Rk545	I0<4>/I1<3>/Q#3	I0<4>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk546	I0<4>/I1<3>/Q#5	I0<4>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk547	I0<4>/I1<3>/Q#4	I0<4>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk548	VDD#325	VDD#326	   68.7306	$metal1_conn
Rk549	VDD#327	VDD#328	   31.6000	$metal1_conn
Rk550	VDD#329	VDD#330	   68.7306	$metal1_conn
Rk551	BLB<36>#3	BLB<36>#1	   75.0000	$metal1_conn
Rk552	I0<4>/I1<3>/QB#4	I0<4>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk553	I0<4>/I1<3>/QB#6	I0<4>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk554	I0<4>/I1<3>/QB#5	I0<4>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk555	WL#147	WL#157	   51.6000	$metal1_conn
Rk556	VSS#223	VSS#4	   19.0550	$metal1_conn
Rk557	VSS#227	VSS#224	   75.1654	$metal1_conn
Rk558	VSS#224	VSS#228	   75.1654	$metal1_conn
Rk559	BLB<37>#1	BLB<37>#2	   81.6000	$metal1_conn
Rk560	I0<4>/I1<6>/QB#3	I0<4>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk561	I0<4>/I1<6>/QB#5	I0<4>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk562	I0<4>/I1<6>/QB#4	I0<4>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk563	VDD#334	VDD#335	   68.7306	$metal1_conn
Rk564	VDD#336	VDD#337	   31.6000	$metal1_conn
Rk565	VDD#338	VDD#339	   68.7306	$metal1_conn
Rk566	BL<37>#1	BL<37>#2	   81.6000	$metal1_conn
Rk567	I0<4>/I1<6>/Q#4	I0<4>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk568	I0<4>/I1<6>/Q#6	I0<4>/I1<6>/Q	    0.1668	$metal1_conn
Rk569	I0<4>/I1<6>/Q#5	I0<4>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk570	WL#151	WL#161	   51.6000	$metal1_conn
Rk571	VSS#231	VSS#4	   19.0550	$metal1_conn
Rk572	VSS#233	VSS#230	   75.1654	$metal1_conn
Rk573	VSS#230	VSS#234	   75.1654	$metal1_conn
Rk574	BL<38>#1	BL<38>#2	   81.6000	$metal1_conn
Rk575	I0<4>/I1<5>/Q#3	I0<4>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk576	I0<4>/I1<5>/Q#5	I0<4>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk577	I0<4>/I1<5>/Q#4	I0<4>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk578	VDD#343	VDD#344	   68.7306	$metal1_conn
Rk579	VDD#345	VDD#346	   31.6000	$metal1_conn
Rk580	VDD#347	VDD#348	   68.7306	$metal1_conn
Rk581	BLB<38>#3	BLB<38>#1	   75.0000	$metal1_conn
Rk582	I0<4>/I1<5>/QB#4	I0<4>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk583	I0<4>/I1<5>/QB#6	I0<4>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk584	I0<4>/I1<5>/QB#5	I0<4>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk585	WL#155	WL#165	   51.6000	$metal1_conn
Rk586	VSS#235	VSS#4	   19.0550	$metal1_conn
Rk587	VSS#239	VSS#236	   75.1654	$metal1_conn
Rk588	VSS#236	VSS#240	   75.1654	$metal1_conn
Rk589	BLB<39>#1	BLB<39>#2	   81.6000	$metal1_conn
Rk590	I0<4>/I1<7>/QB#3	I0<4>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk591	I0<4>/I1<7>/QB#5	I0<4>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk592	I0<4>/I1<7>/QB#4	I0<4>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk593	VDD#352	VDD#353	   68.7306	$metal1_conn
Rk594	VDD#354	VDD#355	   31.6000	$metal1_conn
Rk595	VDD#356	VDD#357	   68.7306	$metal1_conn
Rk596	BL<39>#1	BL<39>#2	   81.6000	$metal1_conn
Rk597	I0<4>/I1<7>/Q#4	I0<4>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk598	I0<4>/I1<7>/Q#6	I0<4>/I1<7>/Q	    0.1668	$metal1_conn
Rk599	I0<4>/I1<7>/Q#5	I0<4>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk600	WL#159	WL#169	   51.6000	$metal1_conn
Rk601	VSS#243	VSS#4	   19.0550	$metal1_conn
Rk602	VSS#245	VSS#242	   75.1654	$metal1_conn
Rk603	VSS#242	VSS#246	   75.1654	$metal1_conn
Rk604	BL<40>#1	BL<40>#2	   81.6000	$metal1_conn
Rk605	I0<5>/I1<0>/Q#3	I0<5>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk606	I0<5>/I1<0>/Q#5	I0<5>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk607	I0<5>/I1<0>/Q#4	I0<5>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk608	VDD#361	VDD#362	   68.7306	$metal1_conn
Rk609	VDD#363	VDD#364	   31.6000	$metal1_conn
Rk610	VDD#365	VDD#366	   68.7306	$metal1_conn
Rk611	BLB<40>#3	BLB<40>#1	   75.0000	$metal1_conn
Rk612	I0<5>/I1<0>/QB#4	I0<5>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk613	I0<5>/I1<0>/QB#6	I0<5>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk614	I0<5>/I1<0>/QB#5	I0<5>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk615	WL#163	WL#173	   51.6000	$metal1_conn
Rk616	VSS#247	VSS#4	   19.0550	$metal1_conn
Rk617	VSS#251	VSS#248	   75.1654	$metal1_conn
Rk618	VSS#248	VSS#252	   75.1654	$metal1_conn
Rk619	BLB<41>#1	BLB<41>#2	   81.6000	$metal1_conn
Rk620	I0<5>/I1<2>/QB#3	I0<5>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk621	I0<5>/I1<2>/QB#5	I0<5>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk622	I0<5>/I1<2>/QB#4	I0<5>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk623	VDD#370	VDD#371	   68.7306	$metal1_conn
Rk624	VDD#372	VDD#373	   31.6000	$metal1_conn
Rk625	VDD#374	VDD#375	   68.7306	$metal1_conn
Rk626	BL<41>#1	BL<41>#2	   81.6000	$metal1_conn
Rk627	I0<5>/I1<2>/Q#4	I0<5>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk628	I0<5>/I1<2>/Q#6	I0<5>/I1<2>/Q	    0.1668	$metal1_conn
Rk629	I0<5>/I1<2>/Q#5	I0<5>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk630	WL#167	WL#177	   51.6000	$metal1_conn
Rk631	VSS#255	VSS#4	   19.0550	$metal1_conn
Rk632	VSS#257	VSS#254	   75.1654	$metal1_conn
Rk633	VSS#254	VSS#258	   75.1654	$metal1_conn
Rk634	BL<42>#1	BL<42>#2	   81.6000	$metal1_conn
Rk635	I0<5>/I1<1>/Q#3	I0<5>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk636	I0<5>/I1<1>/Q#5	I0<5>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk637	I0<5>/I1<1>/Q#4	I0<5>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk638	VDD#379	VDD#380	   68.7306	$metal1_conn
Rk639	VDD#381	VDD#382	   31.6000	$metal1_conn
Rk640	VDD#383	VDD#384	   68.7306	$metal1_conn
Rk641	BLB<42>#3	BLB<42>#1	   75.0000	$metal1_conn
Rk642	I0<5>/I1<1>/QB#4	I0<5>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk643	I0<5>/I1<1>/QB#6	I0<5>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk644	I0<5>/I1<1>/QB#5	I0<5>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk645	WL#171	WL#181	   51.6000	$metal1_conn
Rk646	VSS#259	VSS#4	   19.0550	$metal1_conn
Rk647	VSS#263	VSS#260	   75.1654	$metal1_conn
Rk648	VSS#260	VSS#264	   75.1654	$metal1_conn
Rk649	BLB<43>#1	BLB<43>#2	   81.6000	$metal1_conn
Rk650	I0<5>/I1<4>/QB#3	I0<5>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk651	I0<5>/I1<4>/QB#5	I0<5>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk652	I0<5>/I1<4>/QB#4	I0<5>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk653	VDD#388	VDD#389	   68.7306	$metal1_conn
Rk654	VDD#390	VDD#391	   31.6000	$metal1_conn
Rk655	VDD#392	VDD#393	   68.7306	$metal1_conn
Rk656	BL<43>#1	BL<43>#2	   81.6000	$metal1_conn
Rk657	I0<5>/I1<4>/Q#4	I0<5>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk658	I0<5>/I1<4>/Q#6	I0<5>/I1<4>/Q	    0.1668	$metal1_conn
Rk659	I0<5>/I1<4>/Q#5	I0<5>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk660	WL#175	WL#185	   51.6000	$metal1_conn
Rk661	VSS#267	VSS#4	   19.0550	$metal1_conn
Rk662	VSS#269	VSS#266	   75.1654	$metal1_conn
Rk663	VSS#266	VSS#270	   75.1654	$metal1_conn
Rk664	BL<44>#1	BL<44>#2	   81.6000	$metal1_conn
Rk665	I0<5>/I1<3>/Q#3	I0<5>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk666	I0<5>/I1<3>/Q#5	I0<5>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk667	I0<5>/I1<3>/Q#4	I0<5>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk668	VDD#397	VDD#398	   68.7306	$metal1_conn
Rk669	VDD#399	VDD#400	   31.6000	$metal1_conn
Rk670	VDD#401	VDD#402	   68.7306	$metal1_conn
Rk671	BLB<44>#3	BLB<44>#1	   75.0000	$metal1_conn
Rk672	I0<5>/I1<3>/QB#4	I0<5>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk673	I0<5>/I1<3>/QB#6	I0<5>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk674	I0<5>/I1<3>/QB#5	I0<5>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk675	WL#179	WL#189	   51.6000	$metal1_conn
Rk676	VSS#271	VSS#4	   19.0550	$metal1_conn
Rk677	VSS#275	VSS#272	   75.1654	$metal1_conn
Rk678	VSS#272	VSS#276	   75.1654	$metal1_conn
Rk679	BLB<45>#1	BLB<45>#2	   81.6000	$metal1_conn
Rk680	I0<5>/I1<6>/QB#3	I0<5>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk681	I0<5>/I1<6>/QB#5	I0<5>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk682	I0<5>/I1<6>/QB#4	I0<5>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk683	VDD#406	VDD#407	   68.7306	$metal1_conn
Rk684	VDD#408	VDD#409	   31.6000	$metal1_conn
Rk685	VDD#410	VDD#411	   68.7306	$metal1_conn
Rk686	BL<45>#1	BL<45>#2	   81.6000	$metal1_conn
Rk687	I0<5>/I1<6>/Q#4	I0<5>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk688	I0<5>/I1<6>/Q#6	I0<5>/I1<6>/Q	    0.1668	$metal1_conn
Rk689	I0<5>/I1<6>/Q#5	I0<5>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk690	WL#183	WL#193	   51.6000	$metal1_conn
Rk691	VSS#279	VSS#4	   19.0550	$metal1_conn
Rk692	VSS#281	VSS#278	   75.1654	$metal1_conn
Rk693	VSS#278	VSS#282	   75.1654	$metal1_conn
Rk694	BL<46>#1	BL<46>#2	   81.6000	$metal1_conn
Rk695	I0<5>/I1<5>/Q#3	I0<5>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk696	I0<5>/I1<5>/Q#5	I0<5>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk697	I0<5>/I1<5>/Q#4	I0<5>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk698	VDD#415	VDD#416	   68.7306	$metal1_conn
Rk699	VDD#417	VDD#418	   31.6000	$metal1_conn
Rk700	VDD#419	VDD#420	   68.7306	$metal1_conn
Rk701	BLB<46>#3	BLB<46>#1	   75.0000	$metal1_conn
Rk702	I0<5>/I1<5>/QB#4	I0<5>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk703	I0<5>/I1<5>/QB#6	I0<5>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk704	I0<5>/I1<5>/QB#5	I0<5>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk705	WL#187	WL#197	   51.6000	$metal1_conn
Rk706	VSS#283	VSS#4	   19.0550	$metal1_conn
Rk707	VSS#287	VSS#284	   75.1654	$metal1_conn
Rk708	VSS#284	VSS#288	   75.1654	$metal1_conn
Rk709	BLB<47>#1	BLB<47>#2	   81.6000	$metal1_conn
Rk710	I0<5>/I1<7>/QB#3	I0<5>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk711	I0<5>/I1<7>/QB#5	I0<5>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk712	I0<5>/I1<7>/QB#4	I0<5>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk713	VDD#424	VDD#425	   68.7306	$metal1_conn
Rk714	VDD#426	VDD#427	   31.6000	$metal1_conn
Rk715	VDD#428	VDD#429	   68.7306	$metal1_conn
Rk716	BL<47>#1	BL<47>#2	   81.6000	$metal1_conn
Rk717	I0<5>/I1<7>/Q#4	I0<5>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk718	I0<5>/I1<7>/Q#6	I0<5>/I1<7>/Q	    0.1668	$metal1_conn
Rk719	I0<5>/I1<7>/Q#5	I0<5>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk720	WL#191	WL#201	   51.6000	$metal1_conn
Rk721	VSS#291	VSS#4	   19.0550	$metal1_conn
Rk722	VSS#293	VSS#290	   75.1654	$metal1_conn
Rk723	VSS#290	VSS#294	   75.1654	$metal1_conn
Rk724	BL<48>#1	BL<48>#2	   81.6000	$metal1_conn
Rk725	I0<6>/I1<0>/Q#3	I0<6>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk726	I0<6>/I1<0>/Q#5	I0<6>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk727	I0<6>/I1<0>/Q#4	I0<6>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk728	VDD#433	VDD#434	   68.7306	$metal1_conn
Rk729	VDD#435	VDD#436	   31.6000	$metal1_conn
Rk730	VDD#437	VDD#438	   68.7306	$metal1_conn
Rk731	BLB<48>#3	BLB<48>#1	   75.0000	$metal1_conn
Rk732	I0<6>/I1<0>/QB#4	I0<6>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk733	I0<6>/I1<0>/QB#6	I0<6>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk734	I0<6>/I1<0>/QB#5	I0<6>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk735	WL#195	WL#205	   51.6000	$metal1_conn
Rk736	VSS#295	VSS#4	   19.0550	$metal1_conn
Rk737	VSS#299	VSS#296	   75.1654	$metal1_conn
Rk738	VSS#296	VSS#300	   75.1654	$metal1_conn
Rk739	BLB<49>#1	BLB<49>#2	   81.6000	$metal1_conn
Rk740	I0<6>/I1<2>/QB#3	I0<6>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk741	I0<6>/I1<2>/QB#5	I0<6>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk742	I0<6>/I1<2>/QB#4	I0<6>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk743	VDD#442	VDD#443	   68.7306	$metal1_conn
Rk744	VDD#444	VDD#445	   31.6000	$metal1_conn
Rk745	VDD#446	VDD#447	   68.7306	$metal1_conn
Rk746	BL<49>#1	BL<49>#2	   81.6000	$metal1_conn
Rk747	I0<6>/I1<2>/Q#4	I0<6>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk748	I0<6>/I1<2>/Q#6	I0<6>/I1<2>/Q	    0.1668	$metal1_conn
Rk749	I0<6>/I1<2>/Q#5	I0<6>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk750	WL#199	WL#209	   51.6000	$metal1_conn
Rk751	VSS#303	VSS#4	   19.0550	$metal1_conn
Rk752	VSS#305	VSS#302	   75.1654	$metal1_conn
Rk753	VSS#302	VSS#306	   75.1654	$metal1_conn
Rk754	BL<50>#1	BL<50>#2	   81.6000	$metal1_conn
Rk755	I0<6>/I1<1>/Q#3	I0<6>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk756	I0<6>/I1<1>/Q#5	I0<6>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk757	I0<6>/I1<1>/Q#4	I0<6>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk758	VDD#451	VDD#452	   68.7306	$metal1_conn
Rk759	VDD#453	VDD#454	   31.6000	$metal1_conn
Rk760	VDD#455	VDD#456	   68.7306	$metal1_conn
Rk761	BLB<50>#3	BLB<50>#1	   75.0000	$metal1_conn
Rk762	I0<6>/I1<1>/QB#4	I0<6>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk763	I0<6>/I1<1>/QB#6	I0<6>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk764	I0<6>/I1<1>/QB#5	I0<6>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk765	WL#203	WL#213	   51.6000	$metal1_conn
Rk766	VSS#307	VSS#4	   19.0550	$metal1_conn
Rk767	VSS#311	VSS#308	   75.1654	$metal1_conn
Rk768	VSS#308	VSS#312	   75.1654	$metal1_conn
Rk769	BLB<51>#1	BLB<51>#2	   81.6000	$metal1_conn
Rk770	I0<6>/I1<4>/QB#3	I0<6>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk771	I0<6>/I1<4>/QB#5	I0<6>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk772	I0<6>/I1<4>/QB#4	I0<6>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk773	VDD#460	VDD#461	   68.7306	$metal1_conn
Rk774	VDD#462	VDD#463	   31.6000	$metal1_conn
Rk775	VDD#464	VDD#465	   68.7306	$metal1_conn
Rk776	BL<51>#1	BL<51>#2	   81.6000	$metal1_conn
Rk777	I0<6>/I1<4>/Q#4	I0<6>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk778	I0<6>/I1<4>/Q#6	I0<6>/I1<4>/Q	    0.1668	$metal1_conn
Rk779	I0<6>/I1<4>/Q#5	I0<6>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk780	WL#207	WL#217	   51.6000	$metal1_conn
Rk781	VSS#315	VSS#4	   19.0550	$metal1_conn
Rk782	VSS#317	VSS#314	   75.1654	$metal1_conn
Rk783	VSS#314	VSS#318	   75.1654	$metal1_conn
Rk784	BL<52>#1	BL<52>#2	   81.6000	$metal1_conn
Rk785	I0<6>/I1<3>/Q#3	I0<6>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk786	I0<6>/I1<3>/Q#5	I0<6>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk787	I0<6>/I1<3>/Q#4	I0<6>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk788	VDD#469	VDD#470	   68.7306	$metal1_conn
Rk789	VDD#471	VDD#472	   31.6000	$metal1_conn
Rk790	VDD#473	VDD#474	   68.7306	$metal1_conn
Rk791	BLB<52>#3	BLB<52>#1	   75.0000	$metal1_conn
Rk792	I0<6>/I1<3>/QB#4	I0<6>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk793	I0<6>/I1<3>/QB#6	I0<6>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk794	I0<6>/I1<3>/QB#5	I0<6>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk795	WL#211	WL#221	   51.6000	$metal1_conn
Rk796	VSS#319	VSS#4	   19.0550	$metal1_conn
Rk797	VSS#323	VSS#320	   75.1654	$metal1_conn
Rk798	VSS#320	VSS#324	   75.1654	$metal1_conn
Rk799	BLB<53>#1	BLB<53>#2	   81.6000	$metal1_conn
Rk800	I0<6>/I1<6>/QB#3	I0<6>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk801	I0<6>/I1<6>/QB#5	I0<6>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk802	I0<6>/I1<6>/QB#4	I0<6>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk803	VDD#478	VDD#479	   68.7306	$metal1_conn
Rk804	VDD#480	VDD#481	   31.6000	$metal1_conn
Rk805	VDD#482	VDD#483	   68.7306	$metal1_conn
Rk806	BL<53>#1	BL<53>#2	   81.6000	$metal1_conn
Rk807	I0<6>/I1<6>/Q#4	I0<6>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk808	I0<6>/I1<6>/Q#6	I0<6>/I1<6>/Q	    0.1668	$metal1_conn
Rk809	I0<6>/I1<6>/Q#5	I0<6>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk810	WL#215	WL#225	   51.6000	$metal1_conn
Rk811	VSS#327	VSS#4	   19.0550	$metal1_conn
Rk812	VSS#329	VSS#326	   75.1654	$metal1_conn
Rk813	VSS#326	VSS#330	   75.1654	$metal1_conn
Rk814	BL<54>#1	BL<54>#2	   81.6000	$metal1_conn
Rk815	I0<6>/I1<5>/Q#3	I0<6>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk816	I0<6>/I1<5>/Q#5	I0<6>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk817	I0<6>/I1<5>/Q#4	I0<6>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk818	VDD#487	VDD#488	   68.7306	$metal1_conn
Rk819	VDD#489	VDD#490	   31.6000	$metal1_conn
Rk820	VDD#491	VDD#492	   68.7306	$metal1_conn
Rk821	BLB<54>#3	BLB<54>#1	   75.0000	$metal1_conn
Rk822	I0<6>/I1<5>/QB#4	I0<6>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk823	I0<6>/I1<5>/QB#6	I0<6>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk824	I0<6>/I1<5>/QB#5	I0<6>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk825	WL#219	WL#229	   51.6000	$metal1_conn
Rk826	VSS#331	VSS#4	   19.0550	$metal1_conn
Rk827	VSS#335	VSS#332	   75.1654	$metal1_conn
Rk828	VSS#332	VSS#336	   75.1654	$metal1_conn
Rk829	BLB<55>#1	BLB<55>#2	   81.6000	$metal1_conn
Rk830	I0<6>/I1<7>/QB#3	I0<6>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk831	I0<6>/I1<7>/QB#5	I0<6>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk832	I0<6>/I1<7>/QB#4	I0<6>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk833	VDD#496	VDD#497	   68.7306	$metal1_conn
Rk834	VDD#498	VDD#499	   31.6000	$metal1_conn
Rk835	VDD#500	VDD#501	   68.7306	$metal1_conn
Rk836	BL<55>#1	BL<55>#2	   81.6000	$metal1_conn
Rk837	I0<6>/I1<7>/Q#4	I0<6>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk838	I0<6>/I1<7>/Q#6	I0<6>/I1<7>/Q	    0.1668	$metal1_conn
Rk839	I0<6>/I1<7>/Q#5	I0<6>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk840	WL#223	WL#233	   51.6000	$metal1_conn
Rk841	VSS#339	VSS#4	   19.0550	$metal1_conn
Rk842	VSS#341	VSS#338	   75.1654	$metal1_conn
Rk843	VSS#338	VSS#342	   75.1654	$metal1_conn
Rk844	BL<56>#1	BL<56>#2	   81.6000	$metal1_conn
Rk845	I0<7>/I1<0>/Q#3	I0<7>/I1<0>/Q#5	    0.1668
+ $metal1_conn
Rk846	I0<7>/I1<0>/Q#5	I0<7>/I1<0>/Q#6	   75.2863
+ $metal1_conn
Rk847	I0<7>/I1<0>/Q#4	I0<7>/I1<0>/Q#5	   62.0000
+ $metal1_conn
Rk848	VDD#505	VDD#506	   68.7306	$metal1_conn
Rk849	VDD#507	VDD#508	   31.6000	$metal1_conn
Rk850	VDD#509	VDD#510	   68.7306	$metal1_conn
Rk851	BLB<56>#3	BLB<56>#1	   75.0000	$metal1_conn
Rk852	I0<7>/I1<0>/QB#4	I0<7>/I1<0>/QB#6	   75.2854
+ $metal1_conn
Rk853	I0<7>/I1<0>/QB#6	I0<7>/I1<0>/QB#3	    0.1668
+ $metal1_conn
Rk854	I0<7>/I1<0>/QB#5	I0<7>/I1<0>/QB#6	   62.0000
+ $metal1_conn
Rk855	WL#227	WL#237	   51.6000	$metal1_conn
Rk856	VSS#343	VSS#4	   19.0550	$metal1_conn
Rk857	VSS#347	VSS#344	   75.1654	$metal1_conn
Rk858	VSS#344	VSS#348	   75.1654	$metal1_conn
Rk859	BLB<57>#1	BLB<57>#2	   81.6000	$metal1_conn
Rk860	I0<7>/I1<2>/QB#3	I0<7>/I1<2>/QB#5	    0.1668
+ $metal1_conn
Rk861	I0<7>/I1<2>/QB#5	I0<7>/I1<2>/QB#6	   75.2854
+ $metal1_conn
Rk862	I0<7>/I1<2>/QB#4	I0<7>/I1<2>/QB#5	   62.0000
+ $metal1_conn
Rk863	VDD#514	VDD#515	   68.7306	$metal1_conn
Rk864	VDD#516	VDD#517	   31.6000	$metal1_conn
Rk865	VDD#518	VDD#519	   68.7306	$metal1_conn
Rk866	BL<57>#1	BL<57>#2	   81.6000	$metal1_conn
Rk867	I0<7>/I1<2>/Q#4	I0<7>/I1<2>/Q#6	   75.2863
+ $metal1_conn
Rk868	I0<7>/I1<2>/Q#6	I0<7>/I1<2>/Q	    0.1668	$metal1_conn
Rk869	I0<7>/I1<2>/Q#5	I0<7>/I1<2>/Q#6	   62.0000
+ $metal1_conn
Rk870	WL#231	WL#241	   51.6000	$metal1_conn
Rk871	VSS#351	VSS#4	   19.0550	$metal1_conn
Rk872	VSS#353	VSS#350	   75.1654	$metal1_conn
Rk873	VSS#350	VSS#354	   75.1654	$metal1_conn
Rk874	BL<58>#1	BL<58>#2	   81.6000	$metal1_conn
Rk875	I0<7>/I1<1>/Q#3	I0<7>/I1<1>/Q#5	    0.1668
+ $metal1_conn
Rk876	I0<7>/I1<1>/Q#5	I0<7>/I1<1>/Q#6	   75.2863
+ $metal1_conn
Rk877	I0<7>/I1<1>/Q#4	I0<7>/I1<1>/Q#5	   62.0000
+ $metal1_conn
Rk878	VDD#523	VDD#524	   68.7306	$metal1_conn
Rk879	VDD#525	VDD#526	   31.6000	$metal1_conn
Rk880	VDD#527	VDD#528	   68.7306	$metal1_conn
Rk881	BLB<58>#3	BLB<58>#1	   75.0000	$metal1_conn
Rk882	I0<7>/I1<1>/QB#4	I0<7>/I1<1>/QB#6	   75.2854
+ $metal1_conn
Rk883	I0<7>/I1<1>/QB#6	I0<7>/I1<1>/QB#3	    0.1668
+ $metal1_conn
Rk884	I0<7>/I1<1>/QB#5	I0<7>/I1<1>/QB#6	   62.0000
+ $metal1_conn
Rk885	WL#235	WL#245	   51.6000	$metal1_conn
Rk886	VSS#355	VSS#4	   19.0550	$metal1_conn
Rk887	VSS#359	VSS#356	   75.1654	$metal1_conn
Rk888	VSS#356	VSS#360	   75.1654	$metal1_conn
Rk889	BLB<59>#1	BLB<59>#2	   81.6000	$metal1_conn
Rk890	I0<7>/I1<4>/QB#3	I0<7>/I1<4>/QB#5	    0.1668
+ $metal1_conn
Rk891	I0<7>/I1<4>/QB#5	I0<7>/I1<4>/QB#6	   75.2854
+ $metal1_conn
Rk892	I0<7>/I1<4>/QB#4	I0<7>/I1<4>/QB#5	   62.0000
+ $metal1_conn
Rk893	VDD#532	VDD#533	   68.7306	$metal1_conn
Rk894	VDD#534	VDD#535	   31.6000	$metal1_conn
Rk895	VDD#536	VDD#537	   68.7306	$metal1_conn
Rk896	BL<59>#1	BL<59>#2	   81.6000	$metal1_conn
Rk897	I0<7>/I1<4>/Q#4	I0<7>/I1<4>/Q#6	   75.2863
+ $metal1_conn
Rk898	I0<7>/I1<4>/Q#6	I0<7>/I1<4>/Q	    0.1668	$metal1_conn
Rk899	I0<7>/I1<4>/Q#5	I0<7>/I1<4>/Q#6	   62.0000
+ $metal1_conn
Rk900	WL#239	WL#249	   51.6000	$metal1_conn
Rk901	VSS#363	VSS#4	   19.0550	$metal1_conn
Rk902	VSS#365	VSS#362	   75.1654	$metal1_conn
Rk903	VSS#362	VSS#366	   75.1654	$metal1_conn
Rk904	BL<60>#1	BL<60>#2	   81.6000	$metal1_conn
Rk905	I0<7>/I1<3>/Q#3	I0<7>/I1<3>/Q#5	    0.1668
+ $metal1_conn
Rk906	I0<7>/I1<3>/Q#5	I0<7>/I1<3>/Q#6	   75.2863
+ $metal1_conn
Rk907	I0<7>/I1<3>/Q#4	I0<7>/I1<3>/Q#5	   62.0000
+ $metal1_conn
Rk908	VDD#541	VDD#542	   68.7306	$metal1_conn
Rk909	VDD#543	VDD#544	   31.6000	$metal1_conn
Rk910	VDD#545	VDD#546	   68.7306	$metal1_conn
Rk911	BLB<60>#3	BLB<60>#1	   75.0000	$metal1_conn
Rk912	I0<7>/I1<3>/QB#4	I0<7>/I1<3>/QB#6	   75.2854
+ $metal1_conn
Rk913	I0<7>/I1<3>/QB#6	I0<7>/I1<3>/QB#3	    0.1668
+ $metal1_conn
Rk914	I0<7>/I1<3>/QB#5	I0<7>/I1<3>/QB#6	   62.0000
+ $metal1_conn
Rk915	WL#243	WL#253	   51.6000	$metal1_conn
Rk916	VSS#367	VSS#4	   19.0550	$metal1_conn
Rk917	VSS#371	VSS#368	   75.1654	$metal1_conn
Rk918	VSS#368	VSS#372	   75.1654	$metal1_conn
Rk919	BLB<61>#1	BLB<61>#2	   81.6000	$metal1_conn
Rk920	I0<7>/I1<6>/QB#3	I0<7>/I1<6>/QB#5	    0.1668
+ $metal1_conn
Rk921	I0<7>/I1<6>/QB#5	I0<7>/I1<6>/QB#6	   75.2854
+ $metal1_conn
Rk922	I0<7>/I1<6>/QB#4	I0<7>/I1<6>/QB#5	   62.0000
+ $metal1_conn
Rk923	VDD#550	VDD#551	   68.7306	$metal1_conn
Rk924	VDD#552	VDD#553	   31.6000	$metal1_conn
Rk925	VDD#554	VDD#555	   68.7306	$metal1_conn
Rk926	BL<61>#1	BL<61>#2	   81.6000	$metal1_conn
Rk927	I0<7>/I1<6>/Q#4	I0<7>/I1<6>/Q#6	   75.2863
+ $metal1_conn
Rk928	I0<7>/I1<6>/Q#6	I0<7>/I1<6>/Q	    0.1668	$metal1_conn
Rk929	I0<7>/I1<6>/Q#5	I0<7>/I1<6>/Q#6	   62.0000
+ $metal1_conn
Rk930	WL#247	WL#256	   51.6000	$metal1_conn
Rk931	VSS#373	VSS#4	   19.0550	$metal1_conn
Rk932	VSS#374	VSS#375	   75.1654	$metal1_conn
Rk933	VSS#375	VSS#376	   75.1654	$metal1_conn
Rk934	BL<62>#1	BL<62>#2	   81.6000	$metal1_conn
Rk935	I0<7>/I1<5>/Q#3	I0<7>/I1<5>/Q#5	    0.1668
+ $metal1_conn
Rk936	I0<7>/I1<5>/Q#5	I0<7>/I1<5>/Q#6	   75.2863
+ $metal1_conn
Rk937	I0<7>/I1<5>/Q#4	I0<7>/I1<5>/Q#5	   62.0000
+ $metal1_conn
Rk938	VDD#556	VDD#557	   68.7306	$metal1_conn
Rk939	VDD#558	VDD#559	   31.6000	$metal1_conn
Rk940	VDD#560	VDD#561	   68.7306	$metal1_conn
Rk941	BLB<62>#1	BLB<62>#2	   81.6000	$metal1_conn
Rk942	I0<7>/I1<5>/QB#4	I0<7>/I1<5>/QB#6	   75.2854
+ $metal1_conn
Rk943	I0<7>/I1<5>/QB#6	I0<7>/I1<5>/QB#3	    0.1668
+ $metal1_conn
Rk944	I0<7>/I1<5>/QB#5	I0<7>/I1<5>/QB#6	   62.0000
+ $metal1_conn
Rk945	WL#251	WL#257	   51.6000	$metal1_conn
Rk946	VSS#377	VSS#4	   19.0550	$metal1_conn
Rk947	VSS#378	VSS#379	   75.1654	$metal1_conn
Rk948	VSS#379	VSS#380	   75.1654	$metal1_conn
Rk949	BLB<63>#1	BLB<63>#2	   81.6000	$metal1_conn
Rk950	I0<7>/I1<7>/QB#3	I0<7>/I1<7>/QB#5	    0.1668
+ $metal1_conn
Rk951	I0<7>/I1<7>/QB#5	I0<7>/I1<7>/QB#6	   75.2854
+ $metal1_conn
Rk952	I0<7>/I1<7>/QB#4	I0<7>/I1<7>/QB#5	   62.0000
+ $metal1_conn
Rk953	VDD#562	VDD#563	   68.7306	$metal1_conn
Rk954	VDD#564	VDD#565	   31.6000	$metal1_conn
Rk955	VDD#566	VDD#567	   68.7306	$metal1_conn
Rk956	BL<63>#1	BL<63>#2	   81.6000	$metal1_conn
Rk957	I0<7>/I1<7>/Q#4	I0<7>/I1<7>/Q#6	   75.2863
+ $metal1_conn
Rk958	I0<7>/I1<7>/Q#6	I0<7>/I1<7>/Q	    0.1668	$metal1_conn
Rk959	I0<7>/I1<7>/Q#5	I0<7>/I1<7>/Q#6	   62.0000
+ $metal1_conn
Rk960	WL#255	WL#258	    6.6000	$metal1_conn
Rk961	VSS#381	VSS#4	   27.3718	$metal1_conn
Rk962	VSS#382	VSS#383	   81.7654	$metal1_conn
Rj1	VSS#1	VSS#2	   13.2000	$metal2_conn
Rj2	BL<0>#2	BL<0>#3	    6.6000	$metal2_conn
Rj3	VDD#7	VDD#6	    6.6000	$metal2_conn
Rj4	VDD#1	VDD#8	    6.6000	$metal2_conn
Rj5	BLB<0>#1	BLB<0>#2	   13.2000	$metal2_conn
Rj6	VSS#8	VSS#9	   13.2000	$metal2_conn
Rj7	BLB<1>#3	BLB<1>#2	    6.6000	$metal2_conn
Rj8	VDD#10	VDD#16	    6.6000	$metal2_conn
Rj9	VDD#17	VDD#15	    6.6000	$metal2_conn
Rj10	BL<1>#3	BL<1>#2	    6.6000	$metal2_conn
Rj11	VSS#13	VSS#14	   13.2000	$metal2_conn
Rj12	BL<2>#2	BL<2>#3	    6.6000	$metal2_conn
Rj13	VDD#25	VDD#24	    6.6000	$metal2_conn
Rj14	VDD#19	VDD#26	    6.6000	$metal2_conn
Rj15	BLB<2>#1	BLB<2>#2	   13.2000	$metal2_conn
Rj16	VSS#20	VSS#21	   13.2000	$metal2_conn
Rj17	BLB<3>#3	BLB<3>#2	    6.6000	$metal2_conn
Rj18	VDD#28	VDD#34	    6.6000	$metal2_conn
Rj19	VDD#35	VDD#33	    6.6000	$metal2_conn
Rj20	BL<3>#3	BL<3>#2	    6.6000	$metal2_conn
Rj21	VSS#25	VSS#26	   13.2000	$metal2_conn
Rj22	BL<4>#2	BL<4>#3	    6.6000	$metal2_conn
Rj23	VDD#43	VDD#42	    6.6000	$metal2_conn
Rj24	VDD#37	VDD#44	    6.6000	$metal2_conn
Rj25	BLB<4>#1	BLB<4>#2	   13.2000	$metal2_conn
Rj26	VSS#32	VSS#33	   13.2000	$metal2_conn
Rj27	BLB<5>#3	BLB<5>#2	    6.6000	$metal2_conn
Rj28	VDD#46	VDD#52	    6.6000	$metal2_conn
Rj29	VDD#53	VDD#51	    6.6000	$metal2_conn
Rj30	BL<5>#3	BL<5>#2	    6.6000	$metal2_conn
Rj31	VSS#37	VSS#38	   13.2000	$metal2_conn
Rj32	BL<6>#2	BL<6>#3	    6.6000	$metal2_conn
Rj33	VDD#61	VDD#60	    6.6000	$metal2_conn
Rj34	VDD#55	VDD#62	    6.6000	$metal2_conn
Rj35	BLB<6>#1	BLB<6>#2	   13.2000	$metal2_conn
Rj36	VSS#44	VSS#45	   13.2000	$metal2_conn
Rj37	BLB<7>#3	BLB<7>#2	    6.6000	$metal2_conn
Rj38	VDD#64	VDD#70	    6.6000	$metal2_conn
Rj39	VDD#71	VDD#69	    6.6000	$metal2_conn
Rj40	BL<7>#3	BL<7>#2	    6.6000	$metal2_conn
Rj41	VSS#49	VSS#50	   13.2000	$metal2_conn
Rj42	BL<8>#2	BL<8>#3	    6.6000	$metal2_conn
Rj43	VDD#79	VDD#78	    6.6000	$metal2_conn
Rj44	VDD#73	VDD#80	    6.6000	$metal2_conn
Rj45	BLB<8>#1	BLB<8>#2	   13.2000	$metal2_conn
Rj46	VSS#56	VSS#57	   13.2000	$metal2_conn
Rj47	BLB<9>#3	BLB<9>#2	    6.6000	$metal2_conn
Rj48	VDD#82	VDD#88	    6.6000	$metal2_conn
Rj49	VDD#89	VDD#87	    6.6000	$metal2_conn
Rj50	BL<9>#3	BL<9>#2	    6.6000	$metal2_conn
Rj51	VSS#61	VSS#62	   13.2000	$metal2_conn
Rj52	BL<10>#2	BL<10>#3	    6.6000	$metal2_conn
Rj53	VDD#97	VDD#96	    6.6000	$metal2_conn
Rj54	VDD#91	VDD#98	    6.6000	$metal2_conn
Rj55	BLB<10>#1	BLB<10>#2	   13.2000	$metal2_conn
Rj56	VSS#68	VSS#69	   13.2000	$metal2_conn
Rj57	BLB<11>#3	BLB<11>#2	    6.6000	$metal2_conn
Rj58	VDD#100	VDD#106	    6.6000	$metal2_conn
Rj59	VDD#107	VDD#105	    6.6000	$metal2_conn
Rj60	BL<11>#3	BL<11>#2	    6.6000	$metal2_conn
Rj61	VSS#73	VSS#74	   13.2000	$metal2_conn
Rj62	BL<12>#2	BL<12>#3	    6.6000	$metal2_conn
Rj63	VDD#115	VDD#114	    6.6000	$metal2_conn
Rj64	VDD#109	VDD#116	    6.6000	$metal2_conn
Rj65	BLB<12>#1	BLB<12>#2	   13.2000	$metal2_conn
Rj66	VSS#80	VSS#81	   13.2000	$metal2_conn
Rj67	BLB<13>#3	BLB<13>#2	    6.6000	$metal2_conn
Rj68	VDD#118	VDD#124	    6.6000	$metal2_conn
Rj69	VDD#125	VDD#123	    6.6000	$metal2_conn
Rj70	BL<13>#3	BL<13>#2	    6.6000	$metal2_conn
Rj71	VSS#85	VSS#86	   13.2000	$metal2_conn
Rj72	BL<14>#2	BL<14>#3	    6.6000	$metal2_conn
Rj73	VDD#133	VDD#132	    6.6000	$metal2_conn
Rj74	VDD#127	VDD#134	    6.6000	$metal2_conn
Rj75	BLB<14>#1	BLB<14>#2	   13.2000	$metal2_conn
Rj76	VSS#92	VSS#93	   13.2000	$metal2_conn
Rj77	BLB<15>#3	BLB<15>#2	    6.6000	$metal2_conn
Rj78	VDD#136	VDD#142	    6.6000	$metal2_conn
Rj79	VDD#143	VDD#141	    6.6000	$metal2_conn
Rj80	BL<15>#3	BL<15>#2	    6.6000	$metal2_conn
Rj81	VSS#97	VSS#98	   13.2000	$metal2_conn
Rj82	BL<16>#2	BL<16>#3	    6.6000	$metal2_conn
Rj83	VDD#151	VDD#150	    6.6000	$metal2_conn
Rj84	VDD#145	VDD#152	    6.6000	$metal2_conn
Rj85	BLB<16>#1	BLB<16>#2	   13.2000	$metal2_conn
Rj86	VSS#104	VSS#105	   13.2000	$metal2_conn
Rj87	BLB<17>#3	BLB<17>#2	    6.6000	$metal2_conn
Rj88	VDD#154	VDD#160	    6.6000	$metal2_conn
Rj89	VDD#161	VDD#159	    6.6000	$metal2_conn
Rj90	BL<17>#3	BL<17>#2	    6.6000	$metal2_conn
Rj91	VSS#109	VSS#110	   13.2000	$metal2_conn
Rj92	BL<18>#2	BL<18>#3	    6.6000	$metal2_conn
Rj93	VDD#169	VDD#168	    6.6000	$metal2_conn
Rj94	VDD#163	VDD#170	    6.6000	$metal2_conn
Rj95	BLB<18>#1	BLB<18>#2	   13.2000	$metal2_conn
Rj96	VSS#116	VSS#117	   13.2000	$metal2_conn
Rj97	BLB<19>#3	BLB<19>#2	    6.6000	$metal2_conn
Rj98	VDD#172	VDD#178	    6.6000	$metal2_conn
Rj99	VDD#179	VDD#177	    6.6000	$metal2_conn
Rj100	BL<19>#3	BL<19>#2	    6.6000	$metal2_conn
Rj101	VSS#121	VSS#122	   13.2000	$metal2_conn
Rj102	BL<20>#2	BL<20>#3	    6.6000	$metal2_conn
Rj103	VDD#187	VDD#186	    6.6000	$metal2_conn
Rj104	VDD#181	VDD#188	    6.6000	$metal2_conn
Rj105	BLB<20>#1	BLB<20>#2	   13.2000	$metal2_conn
Rj106	VSS#128	VSS#129	   13.2000	$metal2_conn
Rj107	BLB<21>#3	BLB<21>#2	    6.6000	$metal2_conn
Rj108	VDD#190	VDD#196	    6.6000	$metal2_conn
Rj109	VDD#197	VDD#195	    6.6000	$metal2_conn
Rj110	BL<21>#3	BL<21>#2	    6.6000	$metal2_conn
Rj111	VSS#133	VSS#134	   13.2000	$metal2_conn
Rj112	BL<22>#2	BL<22>#3	    6.6000	$metal2_conn
Rj113	VDD#205	VDD#204	    6.6000	$metal2_conn
Rj114	VDD#199	VDD#206	    6.6000	$metal2_conn
Rj115	BLB<22>#1	BLB<22>#2	   13.2000	$metal2_conn
Rj116	VSS#140	VSS#141	   13.2000	$metal2_conn
Rj117	BLB<23>#3	BLB<23>#2	    6.6000	$metal2_conn
Rj118	VDD#208	VDD#214	    6.6000	$metal2_conn
Rj119	VDD#215	VDD#213	    6.6000	$metal2_conn
Rj120	BL<23>#3	BL<23>#2	    6.6000	$metal2_conn
Rj121	VSS#145	VSS#146	   13.2000	$metal2_conn
Rj122	BL<24>#2	BL<24>#3	    6.6000	$metal2_conn
Rj123	VDD#223	VDD#222	    6.6000	$metal2_conn
Rj124	VDD#217	VDD#224	    6.6000	$metal2_conn
Rj125	BLB<24>#1	BLB<24>#2	   13.2000	$metal2_conn
Rj126	VSS#152	VSS#153	   13.2000	$metal2_conn
Rj127	BLB<25>#3	BLB<25>#2	    6.6000	$metal2_conn
Rj128	VDD#226	VDD#232	    6.6000	$metal2_conn
Rj129	VDD#233	VDD#231	    6.6000	$metal2_conn
Rj130	BL<25>#3	BL<25>#2	    6.6000	$metal2_conn
Rj131	VSS#157	VSS#158	   13.2000	$metal2_conn
Rj132	BL<26>#2	BL<26>#3	    6.6000	$metal2_conn
Rj133	VDD#241	VDD#240	    6.6000	$metal2_conn
Rj134	VDD#235	VDD#242	    6.6000	$metal2_conn
Rj135	BLB<26>#1	BLB<26>#2	   13.2000	$metal2_conn
Rj136	VSS#164	VSS#165	   13.2000	$metal2_conn
Rj137	BLB<27>#3	BLB<27>#2	    6.6000	$metal2_conn
Rj138	VDD#244	VDD#250	    6.6000	$metal2_conn
Rj139	VDD#251	VDD#249	    6.6000	$metal2_conn
Rj140	BL<27>#3	BL<27>#2	    6.6000	$metal2_conn
Rj141	VSS#169	VSS#170	   13.2000	$metal2_conn
Rj142	BL<28>#2	BL<28>#3	    6.6000	$metal2_conn
Rj143	VDD#259	VDD#258	    6.6000	$metal2_conn
Rj144	VDD#253	VDD#260	    6.6000	$metal2_conn
Rj145	BLB<28>#1	BLB<28>#2	   13.2000	$metal2_conn
Rj146	VSS#176	VSS#177	   13.2000	$metal2_conn
Rj147	BLB<29>#3	BLB<29>#2	    6.6000	$metal2_conn
Rj148	VDD#262	VDD#268	    6.6000	$metal2_conn
Rj149	VDD#269	VDD#267	    6.6000	$metal2_conn
Rj150	BL<29>#3	BL<29>#2	    6.6000	$metal2_conn
Rj151	VSS#181	VSS#182	   13.2000	$metal2_conn
Rj152	BL<30>#2	BL<30>#3	    6.6000	$metal2_conn
Rj153	VDD#277	VDD#276	    6.6000	$metal2_conn
Rj154	VDD#271	VDD#278	    6.6000	$metal2_conn
Rj155	BLB<30>#1	BLB<30>#2	   13.2000	$metal2_conn
Rj156	VSS#188	VSS#189	   13.2000	$metal2_conn
Rj157	BLB<31>#3	BLB<31>#2	    6.6000	$metal2_conn
Rj158	VDD#280	VDD#286	    6.6000	$metal2_conn
Rj159	VDD#287	VDD#285	    6.6000	$metal2_conn
Rj160	BL<31>#3	BL<31>#2	    6.6000	$metal2_conn
Rj161	VSS#193	VSS#194	   13.2000	$metal2_conn
Rj162	BL<32>#2	BL<32>#3	    6.6000	$metal2_conn
Rj163	VDD#295	VDD#294	    6.6000	$metal2_conn
Rj164	VDD#289	VDD#296	    6.6000	$metal2_conn
Rj165	BLB<32>#1	BLB<32>#2	   13.2000	$metal2_conn
Rj166	VSS#200	VSS#201	   13.2000	$metal2_conn
Rj167	BLB<33>#3	BLB<33>#2	    6.6000	$metal2_conn
Rj168	VDD#298	VDD#304	    6.6000	$metal2_conn
Rj169	VDD#305	VDD#303	    6.6000	$metal2_conn
Rj170	BL<33>#3	BL<33>#2	    6.6000	$metal2_conn
Rj171	VSS#205	VSS#206	   13.2000	$metal2_conn
Rj172	BL<34>#2	BL<34>#3	    6.6000	$metal2_conn
Rj173	VDD#313	VDD#312	    6.6000	$metal2_conn
Rj174	VDD#307	VDD#314	    6.6000	$metal2_conn
Rj175	BLB<34>#1	BLB<34>#2	   13.2000	$metal2_conn
Rj176	VSS#212	VSS#213	   13.2000	$metal2_conn
Rj177	BLB<35>#3	BLB<35>#2	    6.6000	$metal2_conn
Rj178	VDD#316	VDD#322	    6.6000	$metal2_conn
Rj179	VDD#323	VDD#321	    6.6000	$metal2_conn
Rj180	BL<35>#3	BL<35>#2	    6.6000	$metal2_conn
Rj181	VSS#217	VSS#218	   13.2000	$metal2_conn
Rj182	BL<36>#2	BL<36>#3	    6.6000	$metal2_conn
Rj183	VDD#331	VDD#330	    6.6000	$metal2_conn
Rj184	VDD#325	VDD#332	    6.6000	$metal2_conn
Rj185	BLB<36>#1	BLB<36>#2	   13.2000	$metal2_conn
Rj186	VSS#224	VSS#225	   13.2000	$metal2_conn
Rj187	BLB<37>#3	BLB<37>#2	    6.6000	$metal2_conn
Rj188	VDD#334	VDD#340	    6.6000	$metal2_conn
Rj189	VDD#341	VDD#339	    6.6000	$metal2_conn
Rj190	BL<37>#3	BL<37>#2	    6.6000	$metal2_conn
Rj191	VSS#229	VSS#230	   13.2000	$metal2_conn
Rj192	BL<38>#2	BL<38>#3	    6.6000	$metal2_conn
Rj193	VDD#349	VDD#348	    6.6000	$metal2_conn
Rj194	VDD#343	VDD#350	    6.6000	$metal2_conn
Rj195	BLB<38>#1	BLB<38>#2	   13.2000	$metal2_conn
Rj196	VSS#236	VSS#237	   13.2000	$metal2_conn
Rj197	BLB<39>#3	BLB<39>#2	    6.6000	$metal2_conn
Rj198	VDD#352	VDD#358	    6.6000	$metal2_conn
Rj199	VDD#359	VDD#357	    6.6000	$metal2_conn
Rj200	BL<39>#3	BL<39>#2	    6.6000	$metal2_conn
Rj201	VSS#241	VSS#242	   13.2000	$metal2_conn
Rj202	BL<40>#2	BL<40>#3	    6.6000	$metal2_conn
Rj203	VDD#367	VDD#366	    6.6000	$metal2_conn
Rj204	VDD#361	VDD#368	    6.6000	$metal2_conn
Rj205	BLB<40>#1	BLB<40>#2	   13.2000	$metal2_conn
Rj206	VSS#248	VSS#249	   13.2000	$metal2_conn
Rj207	BLB<41>#3	BLB<41>#2	    6.6000	$metal2_conn
Rj208	VDD#370	VDD#376	    6.6000	$metal2_conn
Rj209	VDD#377	VDD#375	    6.6000	$metal2_conn
Rj210	BL<41>#3	BL<41>#2	    6.6000	$metal2_conn
Rj211	VSS#253	VSS#254	   13.2000	$metal2_conn
Rj212	BL<42>#2	BL<42>#3	    6.6000	$metal2_conn
Rj213	VDD#385	VDD#384	    6.6000	$metal2_conn
Rj214	VDD#379	VDD#386	    6.6000	$metal2_conn
Rj215	BLB<42>#1	BLB<42>#2	   13.2000	$metal2_conn
Rj216	VSS#260	VSS#261	   13.2000	$metal2_conn
Rj217	BLB<43>#3	BLB<43>#2	    6.6000	$metal2_conn
Rj218	VDD#388	VDD#394	    6.6000	$metal2_conn
Rj219	VDD#395	VDD#393	    6.6000	$metal2_conn
Rj220	BL<43>#3	BL<43>#2	    6.6000	$metal2_conn
Rj221	VSS#265	VSS#266	   13.2000	$metal2_conn
Rj222	BL<44>#2	BL<44>#3	    6.6000	$metal2_conn
Rj223	VDD#403	VDD#402	    6.6000	$metal2_conn
Rj224	VDD#397	VDD#404	    6.6000	$metal2_conn
Rj225	BLB<44>#1	BLB<44>#2	   13.2000	$metal2_conn
Rj226	VSS#272	VSS#273	   13.2000	$metal2_conn
Rj227	BLB<45>#3	BLB<45>#2	    6.6000	$metal2_conn
Rj228	VDD#406	VDD#412	    6.6000	$metal2_conn
Rj229	VDD#413	VDD#411	    6.6000	$metal2_conn
Rj230	BL<45>#3	BL<45>#2	    6.6000	$metal2_conn
Rj231	VSS#277	VSS#278	   13.2000	$metal2_conn
Rj232	BL<46>#2	BL<46>#3	    6.6000	$metal2_conn
Rj233	VDD#421	VDD#420	    6.6000	$metal2_conn
Rj234	VDD#415	VDD#422	    6.6000	$metal2_conn
Rj235	BLB<46>#1	BLB<46>#2	   13.2000	$metal2_conn
Rj236	VSS#284	VSS#285	   13.2000	$metal2_conn
Rj237	BLB<47>#3	BLB<47>#2	    6.6000	$metal2_conn
Rj238	VDD#424	VDD#430	    6.6000	$metal2_conn
Rj239	VDD#431	VDD#429	    6.6000	$metal2_conn
Rj240	BL<47>#3	BL<47>#2	    6.6000	$metal2_conn
Rj241	VSS#289	VSS#290	   13.2000	$metal2_conn
Rj242	BL<48>#2	BL<48>#3	    6.6000	$metal2_conn
Rj243	VDD#439	VDD#438	    6.6000	$metal2_conn
Rj244	VDD#433	VDD#440	    6.6000	$metal2_conn
Rj245	BLB<48>#1	BLB<48>#2	   13.2000	$metal2_conn
Rj246	VSS#296	VSS#297	   13.2000	$metal2_conn
Rj247	BLB<49>#3	BLB<49>#2	    6.6000	$metal2_conn
Rj248	VDD#442	VDD#448	    6.6000	$metal2_conn
Rj249	VDD#449	VDD#447	    6.6000	$metal2_conn
Rj250	BL<49>#3	BL<49>#2	    6.6000	$metal2_conn
Rj251	VSS#301	VSS#302	   13.2000	$metal2_conn
Rj252	BL<50>#2	BL<50>#3	    6.6000	$metal2_conn
Rj253	VDD#457	VDD#456	    6.6000	$metal2_conn
Rj254	VDD#451	VDD#458	    6.6000	$metal2_conn
Rj255	BLB<50>#1	BLB<50>#2	   13.2000	$metal2_conn
Rj256	VSS#308	VSS#309	   13.2000	$metal2_conn
Rj257	BLB<51>#3	BLB<51>#2	    6.6000	$metal2_conn
Rj258	VDD#460	VDD#466	    6.6000	$metal2_conn
Rj259	VDD#467	VDD#465	    6.6000	$metal2_conn
Rj260	BL<51>#3	BL<51>#2	    6.6000	$metal2_conn
Rj261	VSS#313	VSS#314	   13.2000	$metal2_conn
Rj262	BL<52>#2	BL<52>#3	    6.6000	$metal2_conn
Rj263	VDD#475	VDD#474	    6.6000	$metal2_conn
Rj264	VDD#469	VDD#476	    6.6000	$metal2_conn
Rj265	BLB<52>#1	BLB<52>#2	   13.2000	$metal2_conn
Rj266	VSS#320	VSS#321	   13.2000	$metal2_conn
Rj267	BLB<53>#3	BLB<53>#2	    6.6000	$metal2_conn
Rj268	VDD#478	VDD#484	    6.6000	$metal2_conn
Rj269	VDD#485	VDD#483	    6.6000	$metal2_conn
Rj270	BL<53>#3	BL<53>#2	    6.6000	$metal2_conn
Rj271	VSS#325	VSS#326	   13.2000	$metal2_conn
Rj272	BL<54>#2	BL<54>#3	    6.6000	$metal2_conn
Rj273	VDD#493	VDD#492	    6.6000	$metal2_conn
Rj274	VDD#487	VDD#494	    6.6000	$metal2_conn
Rj275	BLB<54>#1	BLB<54>#2	   13.2000	$metal2_conn
Rj276	VSS#332	VSS#333	   13.2000	$metal2_conn
Rj277	BLB<55>#3	BLB<55>#2	    6.6000	$metal2_conn
Rj278	VDD#496	VDD#502	    6.6000	$metal2_conn
Rj279	VDD#503	VDD#501	    6.6000	$metal2_conn
Rj280	BL<55>#3	BL<55>#2	    6.6000	$metal2_conn
Rj281	VSS#337	VSS#338	   13.2000	$metal2_conn
Rj282	BL<56>#2	BL<56>#3	    6.6000	$metal2_conn
Rj283	VDD#511	VDD#510	    6.6000	$metal2_conn
Rj284	VDD#505	VDD#512	    6.6000	$metal2_conn
Rj285	BLB<56>#1	BLB<56>#2	   13.2000	$metal2_conn
Rj286	VSS#344	VSS#345	   13.2000	$metal2_conn
Rj287	BLB<57>#3	BLB<57>#2	    6.6000	$metal2_conn
Rj288	VDD#514	VDD#520	    6.6000	$metal2_conn
Rj289	VDD#521	VDD#519	    6.6000	$metal2_conn
Rj290	BL<57>#3	BL<57>#2	    6.6000	$metal2_conn
Rj291	VSS#349	VSS#350	   13.2000	$metal2_conn
Rj292	BL<58>#2	BL<58>#3	    6.6000	$metal2_conn
Rj293	VDD#529	VDD#528	    6.6000	$metal2_conn
Rj294	VDD#523	VDD#530	    6.6000	$metal2_conn
Rj295	BLB<58>#1	BLB<58>#2	   13.2000	$metal2_conn
Rj296	VSS#356	VSS#357	   13.2000	$metal2_conn
Rj297	BLB<59>#3	BLB<59>#2	    6.6000	$metal2_conn
Rj298	VDD#532	VDD#538	    6.6000	$metal2_conn
Rj299	VDD#539	VDD#537	    6.6000	$metal2_conn
Rj300	BL<59>#3	BL<59>#2	    6.6000	$metal2_conn
Rj301	VSS#361	VSS#362	   13.2000	$metal2_conn
Rj302	BL<60>#2	BL<60>#3	    6.6000	$metal2_conn
Rj303	VDD#547	VDD#546	    6.6000	$metal2_conn
Rj304	VDD#541	VDD#548	    6.6000	$metal2_conn
Rj305	BLB<60>#1	BLB<60>#2	   13.2000	$metal2_conn
Rj306	VSS#368	VSS#369	   13.2000	$metal2_conn
Rj307	BLB<61>#3	BLB<61>#2	    6.6000	$metal2_conn
Rj308	VDD#550	VDD#568	    6.6000	$metal2_conn
Rj309	VDD#569	VDD#555	    6.6000	$metal2_conn
Rj310	BL<61>#3	BL<61>#2	    6.6000	$metal2_conn
Rj311	VSS#384	VSS#375	   13.2000	$metal2_conn
Rj312	BL<62>#2	BL<62>#3	    6.6000	$metal2_conn
Rj313	VDD#570	VDD#561	    6.6000	$metal2_conn
Rj314	VDD#556	VDD#571	    6.6000	$metal2_conn
Rj315	BLB<62>#2	BLB<62>#3	    6.6000	$metal2_conn
Rj316	VSS#379	VSS#385	   13.2000	$metal2_conn
Rj317	BLB<63>#3	BLB<63>#2	    6.6000	$metal2_conn
Rj318	VDD#562	VDD#572	    6.6000	$metal2_conn
Rj319	VDD#573	VDD#567	    6.6000	$metal2_conn
Rj320	BL<63>#3	BL<63>#2	    6.6000	$metal2_conn
Rj322	VDD#564	VDD#558	    0.9767	$metal2_conn
Rj324	VDD#558	VDD#552	    0.9767	$metal2_conn
Rj326	VDD#552	VDD#543	    0.9767	$metal2_conn
Rj328	VDD#543	VDD#534	    0.9767	$metal2_conn
Rj330	VDD#534	VDD#525	    0.9767	$metal2_conn
Rj332	VDD#525	VDD#516	    0.9767	$metal2_conn
Rj334	VDD#516	VDD#507	    0.9767	$metal2_conn
Rj336	VDD#507	VDD#498	    0.9767	$metal2_conn
Rj338	VDD#498	VDD#489	    0.9767	$metal2_conn
Rj340	VDD#489	VDD#480	    0.9767	$metal2_conn
Rj342	VDD#480	VDD#471	    0.9767	$metal2_conn
Rj344	VDD#471	VDD#462	    0.9767	$metal2_conn
Rj346	VDD#462	VDD#453	    0.9767	$metal2_conn
Rj348	VDD#453	VDD#444	    0.9767	$metal2_conn
Rj350	VDD#444	VDD#435	    0.9767	$metal2_conn
Rj352	VDD#435	VDD#426	    0.9767	$metal2_conn
Rj354	VDD#426	VDD#417	    0.9767	$metal2_conn
Rj356	VDD#417	VDD#408	    0.9767	$metal2_conn
Rj358	VDD#408	VDD#399	    0.9767	$metal2_conn
Rj360	VDD#399	VDD#390	    0.9767	$metal2_conn
Rj362	VDD#390	VDD#381	    0.9767	$metal2_conn
Rj364	VDD#381	VDD#372	    0.9767	$metal2_conn
Rj366	VDD#372	VDD#363	    0.9767	$metal2_conn
Rj368	VDD#363	VDD#354	    0.9767	$metal2_conn
Rj370	VDD#354	VDD#345	    0.9767	$metal2_conn
Rj372	VDD#345	VDD#336	    0.9767	$metal2_conn
Rj374	VDD#336	VDD#327	    0.9767	$metal2_conn
Rj376	VDD#327	VDD#318	    0.9767	$metal2_conn
Rj378	VDD#318	VDD#309	    0.9767	$metal2_conn
Rj380	VDD#309	VDD#300	    0.9767	$metal2_conn
Rj382	VDD#300	VDD#291	    0.9767	$metal2_conn
Rj384	VDD#291	VDD#282	    0.9767	$metal2_conn
Rj386	VDD#282	VDD#273	    0.9767	$metal2_conn
Rj388	VDD#273	VDD#264	    0.9767	$metal2_conn
Rj390	VDD#264	VDD#255	    0.9767	$metal2_conn
Rj392	VDD#255	VDD#246	    0.9767	$metal2_conn
Rj394	VDD#246	VDD#237	    0.9767	$metal2_conn
Rj396	VDD#237	VDD#228	    0.9767	$metal2_conn
Rj398	VDD#228	VDD#219	    0.9767	$metal2_conn
Rj400	VDD#219	VDD#210	    0.9767	$metal2_conn
Rj402	VDD#210	VDD#201	    0.9767	$metal2_conn
Rj404	VDD#201	VDD#192	    0.9767	$metal2_conn
Rj406	VDD#192	VDD#183	    0.9767	$metal2_conn
Rj408	VDD#183	VDD#174	    0.9767	$metal2_conn
Rj410	VDD#174	VDD#165	    0.9767	$metal2_conn
Rj412	VDD#165	VDD#156	    0.9767	$metal2_conn
Rj414	VDD#156	VDD#147	    0.9767	$metal2_conn
Rj416	VDD#147	VDD#138	    0.9767	$metal2_conn
Rj418	VDD#138	VDD#129	    0.9767	$metal2_conn
Rj420	VDD#129	VDD#120	    0.9767	$metal2_conn
Rj422	VDD#120	VDD#111	    0.9767	$metal2_conn
Rj424	VDD#111	VDD#102	    0.9767	$metal2_conn
Rj426	VDD#102	VDD#93	    0.9767	$metal2_conn
Rj428	VDD#93	VDD#84	    0.9767	$metal2_conn
Rj430	VDD#84	VDD#75	    0.9767	$metal2_conn
Rj432	VDD#75	VDD#66	    0.9767	$metal2_conn
Rj434	VDD#66	VDD#57	    0.9767	$metal2_conn
Rj436	VDD#57	VDD#48	    0.9767	$metal2_conn
Rj438	VDD#48	VDD#39	    0.9767	$metal2_conn
Rj440	VDD#39	VDD#30	    0.9767	$metal2_conn
Rj442	VDD#30	VDD#21	    0.9767	$metal2_conn
Rj444	VDD#21	VDD#12	    0.9767	$metal2_conn
Rj446	VDD#12	VDD#3	    0.9767	$metal2_conn
Rj449	VSS#381	VSS#377	    0.9767	$metal2_conn
Rj451	VSS#377	VSS#373	    0.9767	$metal2_conn
Rj453	VSS#373	VSS#367	    0.9767	$metal2_conn
Rj455	VSS#367	VSS#363	    0.9767	$metal2_conn
Rj457	VSS#363	VSS#355	    0.9767	$metal2_conn
Rj459	VSS#355	VSS#351	    0.9767	$metal2_conn
Rj461	VSS#351	VSS#343	    0.9767	$metal2_conn
Rj463	VSS#343	VSS#339	    0.9767	$metal2_conn
Rj465	VSS#339	VSS#331	    0.9767	$metal2_conn
Rj467	VSS#331	VSS#327	    0.9767	$metal2_conn
Rj469	VSS#327	VSS#319	    0.9767	$metal2_conn
Rj471	VSS#319	VSS#315	    0.9767	$metal2_conn
Rj473	VSS#315	VSS#307	    0.9767	$metal2_conn
Rj475	VSS#307	VSS#303	    0.9767	$metal2_conn
Rj477	VSS#303	VSS#295	    0.9767	$metal2_conn
Rj479	VSS#295	VSS#291	    0.9767	$metal2_conn
Rj481	VSS#291	VSS#283	    0.9767	$metal2_conn
Rj483	VSS#283	VSS#279	    0.9767	$metal2_conn
Rj485	VSS#279	VSS#271	    0.9767	$metal2_conn
Rj487	VSS#271	VSS#267	    0.9767	$metal2_conn
Rj489	VSS#267	VSS#259	    0.9767	$metal2_conn
Rj491	VSS#259	VSS#255	    0.9767	$metal2_conn
Rj493	VSS#255	VSS#247	    0.9767	$metal2_conn
Rj495	VSS#247	VSS#243	    0.9767	$metal2_conn
Rj497	VSS#243	VSS#235	    0.9767	$metal2_conn
Rj499	VSS#235	VSS#231	    0.9767	$metal2_conn
Rj501	VSS#231	VSS#223	    0.9767	$metal2_conn
Rj503	VSS#223	VSS#219	    0.9767	$metal2_conn
Rj505	VSS#219	VSS#211	    0.9767	$metal2_conn
Rj507	VSS#211	VSS#207	    0.9767	$metal2_conn
Rj509	VSS#207	VSS#199	    0.9767	$metal2_conn
Rj511	VSS#199	VSS#195	    0.9767	$metal2_conn
Rj513	VSS#195	VSS#187	    0.9767	$metal2_conn
Rj515	VSS#187	VSS#183	    0.9767	$metal2_conn
Rj517	VSS#183	VSS#175	    0.9767	$metal2_conn
Rj519	VSS#175	VSS#171	    0.9767	$metal2_conn
Rj521	VSS#171	VSS#163	    0.9767	$metal2_conn
Rj523	VSS#163	VSS#159	    0.9767	$metal2_conn
Rj525	VSS#159	VSS#151	    0.9767	$metal2_conn
Rj527	VSS#151	VSS#147	    0.9767	$metal2_conn
Rj529	VSS#147	VSS#139	    0.9767	$metal2_conn
Rj531	VSS#139	VSS#135	    0.9767	$metal2_conn
Rj533	VSS#135	VSS#127	    0.9767	$metal2_conn
Rj535	VSS#127	VSS#123	    0.9767	$metal2_conn
Rj537	VSS#123	VSS#115	    0.9767	$metal2_conn
Rj539	VSS#115	VSS#111	    0.9767	$metal2_conn
Rj541	VSS#111	VSS#103	    0.9767	$metal2_conn
Rj543	VSS#103	VSS#99	    0.9767	$metal2_conn
Rj545	VSS#99	VSS#91	    0.9767	$metal2_conn
Rj547	VSS#91	VSS#87	    0.9767	$metal2_conn
Rj549	VSS#87	VSS#79	    0.9767	$metal2_conn
Rj551	VSS#79	VSS#75	    0.9767	$metal2_conn
Rj553	VSS#75	VSS#67	    0.9767	$metal2_conn
Rj555	VSS#67	VSS#63	    0.9767	$metal2_conn
Rj557	VSS#63	VSS#55	    0.9767	$metal2_conn
Rj559	VSS#55	VSS#51	    0.9767	$metal2_conn
Rj561	VSS#51	VSS#43	    0.9767	$metal2_conn
Rj563	VSS#43	VSS#39	    0.9767	$metal2_conn
Rj565	VSS#39	VSS#31	    0.9767	$metal2_conn
Rj567	VSS#31	VSS#27	    0.9767	$metal2_conn
Rj569	VSS#27	VSS#19	    0.9767	$metal2_conn
Rj571	VSS#19	VSS#15	    0.9767	$metal2_conn
Rj573	VSS#15	VSS#7	    0.9767	$metal2_conn
Rj575	VSS#7	VSS#3	    0.9767	$metal2_conn
Rj577	WL#258	WL	5.092e-02	$metal2_conn
Rj578	WL	WL#259	    0.8733	$metal2_conn
Rj579	WL#259	WL#260	    0.8878	$metal2_conn
Rj580	WL#260	WL#261	    0.8878	$metal2_conn
Rj581	WL#261	WL#262	    0.8878	$metal2_conn
Rj582	WL#262	WL#263	    0.8878	$metal2_conn
Rj583	WL#263	WL#264	    0.8878	$metal2_conn
Rj584	WL#264	WL#265	    0.8878	$metal2_conn
Rj585	WL#265	WL#266	    0.8878	$metal2_conn
Rj586	WL#266	WL#267	    0.8878	$metal2_conn
Rj587	WL#267	WL#268	    0.8878	$metal2_conn
Rj588	WL#268	WL#269	    0.8878	$metal2_conn
Rj589	WL#269	WL#270	    0.8878	$metal2_conn
Rj590	WL#270	WL#271	    0.8878	$metal2_conn
Rj591	WL#271	WL#272	    0.8878	$metal2_conn
Rj592	WL#272	WL#273	    0.8878	$metal2_conn
Rj593	WL#273	WL#274	    0.8878	$metal2_conn
Rj594	WL#274	WL#275	    0.8878	$metal2_conn
Rj595	WL#275	WL#276	    0.8878	$metal2_conn
Rj596	WL#276	WL#277	    0.8878	$metal2_conn
Rj597	WL#277	WL#278	    0.8878	$metal2_conn
Rj598	WL#278	WL#279	    0.8878	$metal2_conn
Rj599	WL#279	WL#280	    0.8878	$metal2_conn
Rj600	WL#280	WL#281	    0.8878	$metal2_conn
Rj601	WL#281	WL#282	    0.8878	$metal2_conn
Rj602	WL#282	WL#283	    0.8878	$metal2_conn
Rj603	WL#283	WL#284	    0.8878	$metal2_conn
Rj604	WL#284	WL#285	    0.8878	$metal2_conn
Rj605	WL#285	WL#286	    0.8878	$metal2_conn
Rj606	WL#286	WL#287	    0.8878	$metal2_conn
Rj607	WL#287	WL#288	    0.8878	$metal2_conn
Rj608	WL#288	WL#289	    0.8878	$metal2_conn
Rj609	WL#289	WL#290	    0.8878	$metal2_conn
Rj610	WL#290	WL#291	    0.8878	$metal2_conn
Rj611	WL#291	WL#292	    0.8878	$metal2_conn
Rj612	WL#292	WL#293	    0.8878	$metal2_conn
Rj613	WL#293	WL#294	    0.8878	$metal2_conn
Rj614	WL#294	WL#295	    0.8878	$metal2_conn
Rj615	WL#295	WL#296	    0.8878	$metal2_conn
Rj616	WL#296	WL#297	    0.8878	$metal2_conn
Rj617	WL#297	WL#298	    0.8878	$metal2_conn
Rj618	WL#298	WL#299	    0.8878	$metal2_conn
Rj619	WL#299	WL#300	    0.8878	$metal2_conn
Rj620	WL#300	WL#301	    0.8878	$metal2_conn
Rj621	WL#301	WL#302	    0.8878	$metal2_conn
Rj622	WL#302	WL#303	    0.8878	$metal2_conn
Rj623	WL#303	WL#304	    0.8878	$metal2_conn
Rj624	WL#304	WL#305	    0.8878	$metal2_conn
Rj625	WL#305	WL#306	    0.8878	$metal2_conn
Rj626	WL#306	WL#307	    0.8878	$metal2_conn
Rj627	WL#307	WL#308	    0.8878	$metal2_conn
Rj628	WL#308	WL#309	    0.8878	$metal2_conn
Rj629	WL#309	WL#310	    0.8878	$metal2_conn
Rj630	WL#310	WL#311	    0.8878	$metal2_conn
Rj631	WL#311	WL#312	    0.8878	$metal2_conn
Rj632	WL#312	WL#313	    0.8878	$metal2_conn
Rj633	WL#313	WL#314	    0.8878	$metal2_conn
Rj634	WL#314	WL#315	    0.8878	$metal2_conn
Rj635	WL#315	WL#316	    0.8878	$metal2_conn
Rj636	WL#316	WL#317	    0.8878	$metal2_conn
Rj637	WL#317	WL#318	    0.8878	$metal2_conn
Rj638	WL#318	WL#319	    0.8878	$metal2_conn
Rj639	WL#319	WL#320	    0.8878	$metal2_conn
Rj640	WL#320	WL#321	    0.8878	$metal2_conn
Rj641	WL#321	WL#9	    0.9182	$metal2_conn
Rj642	WL#259	WL#257	3.591e-02	$metal2_conn
Rj643	WL#260	WL#256	3.591e-02	$metal2_conn
Rj644	WL#261	WL#253	3.591e-02	$metal2_conn
Rj645	WL#262	WL#249	3.591e-02	$metal2_conn
Rj646	WL#263	WL#245	3.591e-02	$metal2_conn
Rj647	WL#264	WL#241	3.591e-02	$metal2_conn
Rj648	WL#265	WL#237	3.591e-02	$metal2_conn
Rj649	WL#266	WL#233	3.591e-02	$metal2_conn
Rj650	WL#267	WL#229	3.591e-02	$metal2_conn
Rj651	WL#268	WL#225	3.591e-02	$metal2_conn
Rj652	WL#269	WL#221	3.591e-02	$metal2_conn
Rj653	WL#270	WL#217	3.591e-02	$metal2_conn
Rj654	WL#271	WL#213	3.591e-02	$metal2_conn
Rj655	WL#272	WL#209	3.591e-02	$metal2_conn
Rj656	WL#273	WL#205	3.591e-02	$metal2_conn
Rj657	WL#274	WL#201	3.591e-02	$metal2_conn
Rj658	WL#275	WL#197	3.591e-02	$metal2_conn
Rj659	WL#276	WL#193	3.591e-02	$metal2_conn
Rj660	WL#277	WL#189	3.591e-02	$metal2_conn
Rj661	WL#278	WL#185	3.591e-02	$metal2_conn
Rj662	WL#279	WL#181	3.591e-02	$metal2_conn
Rj663	WL#280	WL#177	3.591e-02	$metal2_conn
Rj664	WL#281	WL#173	3.591e-02	$metal2_conn
Rj665	WL#282	WL#169	3.591e-02	$metal2_conn
Rj666	WL#283	WL#165	3.591e-02	$metal2_conn
Rj667	WL#284	WL#161	3.591e-02	$metal2_conn
Rj668	WL#285	WL#157	3.591e-02	$metal2_conn
Rj669	WL#286	WL#153	3.591e-02	$metal2_conn
Rj670	WL#287	WL#149	3.591e-02	$metal2_conn
Rj671	WL#288	WL#145	3.591e-02	$metal2_conn
Rj672	WL#289	WL#141	3.591e-02	$metal2_conn
Rj673	WL#290	WL#137	3.591e-02	$metal2_conn
Rj674	WL#291	WL#133	3.591e-02	$metal2_conn
Rj675	WL#292	WL#129	3.591e-02	$metal2_conn
Rj676	WL#293	WL#125	3.591e-02	$metal2_conn
Rj677	WL#294	WL#121	3.591e-02	$metal2_conn
Rj678	WL#295	WL#117	3.591e-02	$metal2_conn
Rj679	WL#296	WL#113	3.591e-02	$metal2_conn
Rj680	WL#297	WL#109	3.591e-02	$metal2_conn
Rj681	WL#298	WL#105	3.591e-02	$metal2_conn
Rj682	WL#299	WL#101	3.591e-02	$metal2_conn
Rj683	WL#300	WL#97	3.591e-02	$metal2_conn
Rj684	WL#301	WL#93	3.591e-02	$metal2_conn
Rj685	WL#302	WL#89	3.591e-02	$metal2_conn
Rj686	WL#303	WL#85	3.591e-02	$metal2_conn
Rj687	WL#304	WL#81	3.591e-02	$metal2_conn
Rj688	WL#305	WL#77	3.591e-02	$metal2_conn
Rj689	WL#306	WL#73	3.591e-02	$metal2_conn
Rj690	WL#307	WL#69	3.591e-02	$metal2_conn
Rj691	WL#308	WL#65	3.591e-02	$metal2_conn
Rj692	WL#309	WL#61	3.591e-02	$metal2_conn
Rj693	WL#310	WL#57	3.591e-02	$metal2_conn
Rj694	WL#311	WL#53	3.591e-02	$metal2_conn
Rj695	WL#312	WL#49	3.591e-02	$metal2_conn
Rj696	WL#313	WL#45	3.591e-02	$metal2_conn
Rj697	WL#314	WL#41	3.591e-02	$metal2_conn
Rj698	WL#315	WL#37	3.591e-02	$metal2_conn
Rj699	WL#316	WL#33	3.591e-02	$metal2_conn
Rj700	WL#317	WL#29	3.591e-02	$metal2_conn
Rj701	WL#318	WL#25	3.591e-02	$metal2_conn
Rj702	WL#319	WL#21	3.591e-02	$metal2_conn
Rj703	WL#320	WL#17	3.591e-02	$metal2_conn
Rj704	WL#321	WL#13	3.591e-02	$metal2_conn
Rj705	VSS#389	VSS#382	    6.6000	$metal2_conn
Ri1	VSS#1	VSS#3	    6.8035	$metal3_conn
Ri2	BL<0>	BL<0>#3	    0.2568	$metal3_conn
Ri3	VDD#7	VDD#8	    0.2084	$metal3_conn
Ri4	VDD#8	VDD#3	    6.7371	$metal3_conn
Ri5	BLB<0>	BLB<0>#2	4.192e-02	$metal3_conn
Ri6	VSS#9	VSS#7	    7.0183	$metal3_conn
Ri7	BLB<1>	BLB<1>#3	4.192e-02	$metal3_conn
Ri8	VDD#16	VDD#17	    0.2084	$metal3_conn
Ri9	VDD#17	VDD#12	    6.7371	$metal3_conn
Ri10	BL<1>	BL<1>#3	    0.2568	$metal3_conn
Ri11	VSS#13	VSS#15	    6.8035	$metal3_conn
Ri12	BL<2>	BL<2>#3	    0.2568	$metal3_conn
Ri13	VDD#25	VDD#26	    0.2084	$metal3_conn
Ri14	VDD#26	VDD#21	    6.7371	$metal3_conn
Ri15	BLB<2>	BLB<2>#2	4.192e-02	$metal3_conn
Ri16	VSS#21	VSS#19	    7.0183	$metal3_conn
Ri17	BLB<3>	BLB<3>#3	4.192e-02	$metal3_conn
Ri18	VDD#34	VDD#35	    0.2084	$metal3_conn
Ri19	VDD#35	VDD#30	    6.7371	$metal3_conn
Ri20	BL<3>	BL<3>#3	    0.2568	$metal3_conn
Ri21	VSS#25	VSS#27	    6.8035	$metal3_conn
Ri22	BL<4>	BL<4>#3	    0.2568	$metal3_conn
Ri23	VDD#43	VDD#44	    0.2084	$metal3_conn
Ri24	VDD#44	VDD#39	    6.7371	$metal3_conn
Ri25	BLB<4>	BLB<4>#2	4.192e-02	$metal3_conn
Ri26	VSS#33	VSS#31	    7.0183	$metal3_conn
Ri27	BLB<5>	BLB<5>#3	4.192e-02	$metal3_conn
Ri28	VDD#52	VDD#53	    0.2084	$metal3_conn
Ri29	VDD#53	VDD#48	    6.7371	$metal3_conn
Ri30	BL<5>	BL<5>#3	    0.2568	$metal3_conn
Ri31	VSS#37	VSS#39	    6.8035	$metal3_conn
Ri32	BL<6>	BL<6>#3	    0.2568	$metal3_conn
Ri33	VDD#61	VDD#62	    0.2084	$metal3_conn
Ri34	VDD#62	VDD#57	    6.7371	$metal3_conn
Ri35	BLB<6>	BLB<6>#2	4.192e-02	$metal3_conn
Ri36	VSS#45	VSS#43	    7.0183	$metal3_conn
Ri37	BLB<7>	BLB<7>#3	4.192e-02	$metal3_conn
Ri38	VDD#70	VDD#71	    0.2084	$metal3_conn
Ri39	VDD#71	VDD#66	    6.7371	$metal3_conn
Ri40	BL<7>	BL<7>#3	    0.2568	$metal3_conn
Ri41	VSS#49	VSS#51	    6.8035	$metal3_conn
Ri42	BL<8>	BL<8>#3	    0.2568	$metal3_conn
Ri43	VDD#79	VDD#80	    0.2084	$metal3_conn
Ri44	VDD#80	VDD#75	    6.7371	$metal3_conn
Ri45	BLB<8>	BLB<8>#2	4.192e-02	$metal3_conn
Ri46	VSS#57	VSS#55	    7.0183	$metal3_conn
Ri47	BLB<9>	BLB<9>#3	4.192e-02	$metal3_conn
Ri48	VDD#88	VDD#89	    0.2084	$metal3_conn
Ri49	VDD#89	VDD#84	    6.7371	$metal3_conn
Ri50	BL<9>	BL<9>#3	    0.2568	$metal3_conn
Ri51	VSS#61	VSS#63	    6.8035	$metal3_conn
Ri52	BL<10>	BL<10>#3	    0.2568	$metal3_conn
Ri53	VDD#97	VDD#98	    0.2084	$metal3_conn
Ri54	VDD#98	VDD#93	    6.7371	$metal3_conn
Ri55	BLB<10>	BLB<10>#2	4.192e-02	$metal3_conn
Ri56	VSS#69	VSS#67	    7.0183	$metal3_conn
Ri57	BLB<11>	BLB<11>#3	4.192e-02	$metal3_conn
Ri58	VDD#106	VDD#107	    0.2084	$metal3_conn
Ri59	VDD#107	VDD#102	    6.7371	$metal3_conn
Ri60	BL<11>	BL<11>#3	    0.2568	$metal3_conn
Ri61	VSS#73	VSS#75	    6.8035	$metal3_conn
Ri62	BL<12>	BL<12>#3	    0.2568	$metal3_conn
Ri63	VDD#115	VDD#116	    0.2084	$metal3_conn
Ri64	VDD#116	VDD#111	    6.7371	$metal3_conn
Ri65	BLB<12>	BLB<12>#2	4.192e-02	$metal3_conn
Ri66	VSS#81	VSS#79	    7.0183	$metal3_conn
Ri67	BLB<13>	BLB<13>#3	4.192e-02	$metal3_conn
Ri68	VDD#124	VDD#125	    0.2084	$metal3_conn
Ri69	VDD#125	VDD#120	    6.7371	$metal3_conn
Ri70	BL<13>	BL<13>#3	    0.2568	$metal3_conn
Ri71	VSS#85	VSS#87	    6.8035	$metal3_conn
Ri72	BL<14>	BL<14>#3	    0.2568	$metal3_conn
Ri73	VDD#133	VDD#134	    0.2084	$metal3_conn
Ri74	VDD#134	VDD#129	    6.7371	$metal3_conn
Ri75	BLB<14>	BLB<14>#2	4.192e-02	$metal3_conn
Ri76	VSS#93	VSS#91	    7.0183	$metal3_conn
Ri77	BLB<15>	BLB<15>#3	4.192e-02	$metal3_conn
Ri78	VDD#142	VDD#143	    0.2084	$metal3_conn
Ri79	VDD#143	VDD#138	    6.7371	$metal3_conn
Ri80	BL<15>	BL<15>#3	    0.2568	$metal3_conn
Ri81	VSS#97	VSS#99	    6.8035	$metal3_conn
Ri82	BL<16>	BL<16>#3	    0.2568	$metal3_conn
Ri83	VDD#151	VDD#152	    0.2084	$metal3_conn
Ri84	VDD#152	VDD#147	    6.7371	$metal3_conn
Ri85	BLB<16>	BLB<16>#2	4.192e-02	$metal3_conn
Ri86	VSS#105	VSS#103	    7.0183	$metal3_conn
Ri87	BLB<17>	BLB<17>#3	4.192e-02	$metal3_conn
Ri88	VDD#160	VDD#161	    0.2084	$metal3_conn
Ri89	VDD#161	VDD#156	    6.7371	$metal3_conn
Ri90	BL<17>	BL<17>#3	    0.2568	$metal3_conn
Ri91	VSS#109	VSS#111	    6.8035	$metal3_conn
Ri92	BL<18>	BL<18>#3	    0.2568	$metal3_conn
Ri93	VDD#169	VDD#170	    0.2084	$metal3_conn
Ri94	VDD#170	VDD#165	    6.7371	$metal3_conn
Ri95	BLB<18>	BLB<18>#2	4.192e-02	$metal3_conn
Ri96	VSS#117	VSS#115	    7.0183	$metal3_conn
Ri97	BLB<19>	BLB<19>#3	4.192e-02	$metal3_conn
Ri98	VDD#178	VDD#179	    0.2084	$metal3_conn
Ri99	VDD#179	VDD#174	    6.7371	$metal3_conn
Ri100	BL<19>	BL<19>#3	    0.2568	$metal3_conn
Ri101	VSS#121	VSS#123	    6.8035	$metal3_conn
Ri102	BL<20>	BL<20>#3	    0.2568	$metal3_conn
Ri103	VDD#187	VDD#188	    0.2084	$metal3_conn
Ri104	VDD#188	VDD#183	    6.7371	$metal3_conn
Ri105	BLB<20>	BLB<20>#2	4.192e-02	$metal3_conn
Ri106	VSS#129	VSS#127	    7.0183	$metal3_conn
Ri107	BLB<21>	BLB<21>#3	4.192e-02	$metal3_conn
Ri108	VDD#196	VDD#197	    0.2084	$metal3_conn
Ri109	VDD#197	VDD#192	    6.7371	$metal3_conn
Ri110	BL<21>	BL<21>#3	    0.2568	$metal3_conn
Ri111	VSS#133	VSS#135	    6.8035	$metal3_conn
Ri112	BL<22>	BL<22>#3	    0.2568	$metal3_conn
Ri113	VDD#205	VDD#206	    0.2084	$metal3_conn
Ri114	VDD#206	VDD#201	    6.7371	$metal3_conn
Ri115	BLB<22>	BLB<22>#2	4.192e-02	$metal3_conn
Ri116	VSS#141	VSS#139	    7.0183	$metal3_conn
Ri117	BLB<23>	BLB<23>#3	4.192e-02	$metal3_conn
Ri118	VDD#214	VDD#215	    0.2084	$metal3_conn
Ri119	VDD#215	VDD#210	    6.7371	$metal3_conn
Ri120	BL<23>	BL<23>#3	    0.2568	$metal3_conn
Ri121	VSS#145	VSS#147	    6.8035	$metal3_conn
Ri122	BL<24>	BL<24>#3	    0.2568	$metal3_conn
Ri123	VDD#223	VDD#224	    0.2084	$metal3_conn
Ri124	VDD#224	VDD#219	    6.7371	$metal3_conn
Ri125	BLB<24>	BLB<24>#2	4.192e-02	$metal3_conn
Ri126	VSS#153	VSS#151	    7.0183	$metal3_conn
Ri127	BLB<25>	BLB<25>#3	4.192e-02	$metal3_conn
Ri128	VDD#232	VDD#233	    0.2084	$metal3_conn
Ri129	VDD#233	VDD#228	    6.7371	$metal3_conn
Ri130	BL<25>	BL<25>#3	    0.2568	$metal3_conn
Ri131	VSS#157	VSS#159	    6.8035	$metal3_conn
Ri132	BL<26>	BL<26>#3	    0.2568	$metal3_conn
Ri133	VDD#241	VDD#242	    0.2084	$metal3_conn
Ri134	VDD#242	VDD#237	    6.7371	$metal3_conn
Ri135	BLB<26>	BLB<26>#2	4.192e-02	$metal3_conn
Ri136	VSS#165	VSS#163	    7.0183	$metal3_conn
Ri137	BLB<27>	BLB<27>#3	4.192e-02	$metal3_conn
Ri138	VDD#250	VDD#251	    0.2084	$metal3_conn
Ri139	VDD#251	VDD#246	    6.7371	$metal3_conn
Ri140	BL<27>	BL<27>#3	    0.2568	$metal3_conn
Ri141	VSS#169	VSS#171	    6.8035	$metal3_conn
Ri142	BL<28>	BL<28>#3	    0.2568	$metal3_conn
Ri143	VDD#259	VDD#260	    0.2084	$metal3_conn
Ri144	VDD#260	VDD#255	    6.7371	$metal3_conn
Ri145	BLB<28>	BLB<28>#2	4.192e-02	$metal3_conn
Ri146	VSS#177	VSS#175	    7.0183	$metal3_conn
Ri147	BLB<29>	BLB<29>#3	4.192e-02	$metal3_conn
Ri148	VDD#268	VDD#269	    0.2084	$metal3_conn
Ri149	VDD#269	VDD#264	    6.7371	$metal3_conn
Ri150	BL<29>	BL<29>#3	    0.2568	$metal3_conn
Ri151	VSS#181	VSS#183	    6.8035	$metal3_conn
Ri152	BL<30>	BL<30>#3	    0.2568	$metal3_conn
Ri153	VDD#277	VDD#278	    0.2084	$metal3_conn
Ri154	VDD#278	VDD#273	    6.7371	$metal3_conn
Ri155	BLB<30>	BLB<30>#2	4.192e-02	$metal3_conn
Ri156	VSS#189	VSS#187	    7.0183	$metal3_conn
Ri157	BLB<31>	BLB<31>#3	4.192e-02	$metal3_conn
Ri158	VDD#286	VDD#287	    0.2084	$metal3_conn
Ri159	VDD#287	VDD#282	    6.7371	$metal3_conn
Ri160	BL<31>	BL<31>#3	    0.2568	$metal3_conn
Ri161	VSS#193	VSS#195	    6.8035	$metal3_conn
Ri162	BL<32>	BL<32>#3	    0.2568	$metal3_conn
Ri163	VDD#295	VDD#296	    0.2084	$metal3_conn
Ri164	VDD#296	VDD#291	    6.7371	$metal3_conn
Ri165	BLB<32>	BLB<32>#2	4.192e-02	$metal3_conn
Ri166	VSS#201	VSS#199	    7.0183	$metal3_conn
Ri167	BLB<33>	BLB<33>#3	4.192e-02	$metal3_conn
Ri168	VDD#304	VDD#305	    0.2084	$metal3_conn
Ri169	VDD#305	VDD#300	    6.7371	$metal3_conn
Ri170	BL<33>	BL<33>#3	    0.2568	$metal3_conn
Ri171	VSS#205	VSS#207	    6.8035	$metal3_conn
Ri172	BL<34>	BL<34>#3	    0.2568	$metal3_conn
Ri173	VDD#313	VDD#314	    0.2084	$metal3_conn
Ri174	VDD#314	VDD#309	    6.7371	$metal3_conn
Ri175	BLB<34>	BLB<34>#2	4.192e-02	$metal3_conn
Ri176	VSS#213	VSS#211	    7.0183	$metal3_conn
Ri177	BLB<35>	BLB<35>#3	4.192e-02	$metal3_conn
Ri178	VDD#322	VDD#323	    0.2084	$metal3_conn
Ri179	VDD#323	VDD#318	    6.7371	$metal3_conn
Ri180	BL<35>	BL<35>#3	    0.2568	$metal3_conn
Ri181	VSS#217	VSS#219	    6.8035	$metal3_conn
Ri182	BL<36>	BL<36>#3	    0.2568	$metal3_conn
Ri183	VDD#331	VDD#332	    0.2084	$metal3_conn
Ri184	VDD#332	VDD#327	    6.7371	$metal3_conn
Ri185	BLB<36>	BLB<36>#2	4.192e-02	$metal3_conn
Ri186	VSS#225	VSS#223	    7.0183	$metal3_conn
Ri187	BLB<37>	BLB<37>#3	4.192e-02	$metal3_conn
Ri188	VDD#340	VDD#341	    0.2084	$metal3_conn
Ri189	VDD#341	VDD#336	    6.7371	$metal3_conn
Ri190	BL<37>	BL<37>#3	    0.2568	$metal3_conn
Ri191	VSS#229	VSS#231	    6.8035	$metal3_conn
Ri192	BL<38>	BL<38>#3	    0.2568	$metal3_conn
Ri193	VDD#349	VDD#350	    0.2084	$metal3_conn
Ri194	VDD#350	VDD#345	    6.7371	$metal3_conn
Ri195	BLB<38>	BLB<38>#2	4.192e-02	$metal3_conn
Ri196	VSS#237	VSS#235	    7.0183	$metal3_conn
Ri197	BLB<39>	BLB<39>#3	4.192e-02	$metal3_conn
Ri198	VDD#358	VDD#359	    0.2084	$metal3_conn
Ri199	VDD#359	VDD#354	    6.7371	$metal3_conn
Ri200	BL<39>	BL<39>#3	    0.2568	$metal3_conn
Ri201	VSS#241	VSS#243	    6.8035	$metal3_conn
Ri202	BL<40>	BL<40>#3	    0.2568	$metal3_conn
Ri203	VDD#367	VDD#368	    0.2084	$metal3_conn
Ri204	VDD#368	VDD#363	    6.7371	$metal3_conn
Ri205	BLB<40>	BLB<40>#2	4.192e-02	$metal3_conn
Ri206	VSS#249	VSS#247	    7.0183	$metal3_conn
Ri207	BLB<41>	BLB<41>#3	4.192e-02	$metal3_conn
Ri208	VDD#376	VDD#377	    0.2084	$metal3_conn
Ri209	VDD#377	VDD#372	    6.7371	$metal3_conn
Ri210	BL<41>	BL<41>#3	    0.2568	$metal3_conn
Ri211	VSS#253	VSS#255	    6.8035	$metal3_conn
Ri212	BL<42>	BL<42>#3	    0.2568	$metal3_conn
Ri213	VDD#385	VDD#386	    0.2084	$metal3_conn
Ri214	VDD#386	VDD#381	    6.7371	$metal3_conn
Ri215	BLB<42>	BLB<42>#2	4.192e-02	$metal3_conn
Ri216	VSS#261	VSS#259	    7.0183	$metal3_conn
Ri217	BLB<43>	BLB<43>#3	4.192e-02	$metal3_conn
Ri218	VDD#394	VDD#395	    0.2084	$metal3_conn
Ri219	VDD#395	VDD#390	    6.7371	$metal3_conn
Ri220	BL<43>	BL<43>#3	    0.2568	$metal3_conn
Ri221	VSS#265	VSS#267	    6.8035	$metal3_conn
Ri222	BL<44>	BL<44>#3	    0.2568	$metal3_conn
Ri223	VDD#403	VDD#404	    0.2084	$metal3_conn
Ri224	VDD#404	VDD#399	    6.7371	$metal3_conn
Ri225	BLB<44>	BLB<44>#2	4.192e-02	$metal3_conn
Ri226	VSS#273	VSS#271	    7.0183	$metal3_conn
Ri227	BLB<45>	BLB<45>#3	4.192e-02	$metal3_conn
Ri228	VDD#412	VDD#413	    0.2084	$metal3_conn
Ri229	VDD#413	VDD#408	    6.7371	$metal3_conn
Ri230	BL<45>	BL<45>#3	    0.2568	$metal3_conn
Ri231	VSS#277	VSS#279	    6.8035	$metal3_conn
Ri232	BL<46>	BL<46>#3	    0.2568	$metal3_conn
Ri233	VDD#421	VDD#422	    0.2084	$metal3_conn
Ri234	VDD#422	VDD#417	    6.7371	$metal3_conn
Ri235	BLB<46>	BLB<46>#2	4.192e-02	$metal3_conn
Ri236	VSS#285	VSS#283	    7.0183	$metal3_conn
Ri237	BLB<47>	BLB<47>#3	4.192e-02	$metal3_conn
Ri238	VDD#430	VDD#431	    0.2084	$metal3_conn
Ri239	VDD#431	VDD#426	    6.7371	$metal3_conn
Ri240	BL<47>	BL<47>#3	    0.2568	$metal3_conn
Ri241	VSS#289	VSS#291	    6.8035	$metal3_conn
Ri242	BL<48>	BL<48>#3	    0.2568	$metal3_conn
Ri243	VDD#439	VDD#440	    0.2084	$metal3_conn
Ri244	VDD#440	VDD#435	    6.7371	$metal3_conn
Ri245	BLB<48>	BLB<48>#2	4.192e-02	$metal3_conn
Ri246	VSS#297	VSS#295	    7.0183	$metal3_conn
Ri247	BLB<49>	BLB<49>#3	4.192e-02	$metal3_conn
Ri248	VDD#448	VDD#449	    0.2084	$metal3_conn
Ri249	VDD#449	VDD#444	    6.7371	$metal3_conn
Ri250	BL<49>	BL<49>#3	    0.2568	$metal3_conn
Ri251	VSS#301	VSS#303	    6.8035	$metal3_conn
Ri252	BL<50>	BL<50>#3	    0.2568	$metal3_conn
Ri253	VDD#457	VDD#458	    0.2084	$metal3_conn
Ri254	VDD#458	VDD#453	    6.7371	$metal3_conn
Ri255	BLB<50>	BLB<50>#2	4.192e-02	$metal3_conn
Ri256	VSS#309	VSS#307	    7.0183	$metal3_conn
Ri257	BLB<51>	BLB<51>#3	4.192e-02	$metal3_conn
Ri258	VDD#466	VDD#467	    0.2084	$metal3_conn
Ri259	VDD#467	VDD#462	    6.7371	$metal3_conn
Ri260	BL<51>	BL<51>#3	    0.2568	$metal3_conn
Ri261	VSS#313	VSS#315	    6.8035	$metal3_conn
Ri262	BL<52>	BL<52>#3	    0.2568	$metal3_conn
Ri263	VDD#475	VDD#476	    0.2084	$metal3_conn
Ri264	VDD#476	VDD#471	    6.7371	$metal3_conn
Ri265	BLB<52>	BLB<52>#2	4.192e-02	$metal3_conn
Ri266	VSS#321	VSS#319	    7.0183	$metal3_conn
Ri267	BLB<53>	BLB<53>#3	4.192e-02	$metal3_conn
Ri268	VDD#484	VDD#485	    0.2084	$metal3_conn
Ri269	VDD#485	VDD#480	    6.7371	$metal3_conn
Ri270	BL<53>	BL<53>#3	    0.2568	$metal3_conn
Ri271	VSS#325	VSS#327	    6.8035	$metal3_conn
Ri272	BL<54>	BL<54>#3	    0.2568	$metal3_conn
Ri273	VDD#493	VDD#494	    0.2084	$metal3_conn
Ri274	VDD#494	VDD#489	    6.7371	$metal3_conn
Ri275	BLB<54>	BLB<54>#2	4.192e-02	$metal3_conn
Ri276	VSS#333	VSS#331	    7.0183	$metal3_conn
Ri277	BLB<55>	BLB<55>#3	4.192e-02	$metal3_conn
Ri278	VDD#502	VDD#503	    0.2084	$metal3_conn
Ri279	VDD#503	VDD#498	    6.7371	$metal3_conn
Ri280	BL<55>	BL<55>#3	    0.2568	$metal3_conn
Ri281	VSS#337	VSS#339	    6.8035	$metal3_conn
Ri282	BL<56>	BL<56>#3	    0.2568	$metal3_conn
Ri283	VDD#511	VDD#512	    0.2084	$metal3_conn
Ri284	VDD#512	VDD#507	    6.7371	$metal3_conn
Ri285	BLB<56>	BLB<56>#2	4.192e-02	$metal3_conn
Ri286	VSS#345	VSS#343	    7.0183	$metal3_conn
Ri287	BLB<57>	BLB<57>#3	4.192e-02	$metal3_conn
Ri288	VDD#520	VDD#521	    0.2084	$metal3_conn
Ri289	VDD#521	VDD#516	    6.7371	$metal3_conn
Ri290	BL<57>	BL<57>#3	    0.2568	$metal3_conn
Ri291	VSS#349	VSS#351	    6.8035	$metal3_conn
Ri292	BL<58>	BL<58>#3	    0.2568	$metal3_conn
Ri293	VDD#529	VDD#530	    0.2084	$metal3_conn
Ri294	VDD#530	VDD#525	    6.7371	$metal3_conn
Ri295	BLB<58>	BLB<58>#2	4.192e-02	$metal3_conn
Ri296	VSS#357	VSS#355	    7.0183	$metal3_conn
Ri297	BLB<59>	BLB<59>#3	4.192e-02	$metal3_conn
Ri298	VDD#538	VDD#539	    0.2084	$metal3_conn
Ri299	VDD#539	VDD#534	    6.7371	$metal3_conn
Ri300	BL<59>	BL<59>#3	    0.2568	$metal3_conn
Ri301	VSS#361	VSS#363	    6.8035	$metal3_conn
Ri302	BL<60>	BL<60>#3	    0.2568	$metal3_conn
Ri303	VDD#547	VDD#548	    0.2084	$metal3_conn
Ri304	VDD#548	VDD#543	    6.7371	$metal3_conn
Ri305	BLB<60>	BLB<60>#2	4.192e-02	$metal3_conn
Ri306	VSS#369	VSS#367	    7.0183	$metal3_conn
Ri307	BLB<61>	BLB<61>#3	4.192e-02	$metal3_conn
Ri308	VDD#568	VDD#569	    0.2084	$metal3_conn
Ri309	VDD#569	VDD#552	    6.7371	$metal3_conn
Ri310	BL<61>	BL<61>#3	    0.2568	$metal3_conn
Ri311	VSS#384	VSS#373	    6.8035	$metal3_conn
Ri312	BL<62>	BL<62>#3	    0.2568	$metal3_conn
Ri313	VDD#570	VDD#571	    0.2084	$metal3_conn
Ri314	VDD#571	VDD#558	    6.7371	$metal3_conn
Ri315	BLB<62>	BLB<62>#3	4.192e-02	$metal3_conn
Ri316	VSS	VSS#377	    6.7615	$metal3_conn
Ri317	VSS	VSS#385	    0.2568	$metal3_conn
Ri318	BLB<63>	BLB<63>#3	4.192e-02	$metal3_conn
Ri319	VDD	VDD#564	    6.6977	$metal3_conn
Ri320	VDD	VDD#573	3.949e-02	$metal3_conn
Ri321	VDD#573	VDD#572	    0.2084	$metal3_conn
Ri322	BL<63>	BL<63>#3	    0.2568	$metal3_conn
Ri323	VSS#389	VSS#381	    6.8035	$metal3_conn
*
*       CAPACITOR CARDS
*
*
C1	VDD	VSS	7.81019e-18	$cmodel
C2	WL	VSS	1.33376e-16	$cmodel
C3	BL<0>	VSS	4.00738e-17	$cmodel
C4	BL<10>	VSS	4.00324e-17	$cmodel
C5	BL<11>	VSS	4.00835e-17	$cmodel
C6	BL<12>	VSS	4.00324e-17	$cmodel
C7	BL<13>	VSS	4.00835e-17	$cmodel
C8	BL<14>	VSS	4.00324e-17	$cmodel
C9	BL<15>	VSS	4.00835e-17	$cmodel
C10	BL<16>	VSS	4.00324e-17	$cmodel
C11	BL<17>	VSS	4.00835e-17	$cmodel
C12	BL<18>	VSS	4.00324e-17	$cmodel
C13	BL<19>	VSS	4.00835e-17	$cmodel
C14	BL<1>	VSS	4.00835e-17	$cmodel
C15	BL<20>	VSS	4.00324e-17	$cmodel
C16	BL<21>	VSS	4.00835e-17	$cmodel
C17	BL<22>	VSS	4.00324e-17	$cmodel
C18	BL<23>	VSS	4.00835e-17	$cmodel
C19	BL<24>	VSS	4.00324e-17	$cmodel
C20	BL<25>	VSS	4.00835e-17	$cmodel
C21	BL<26>	VSS	4.00324e-17	$cmodel
C22	BL<27>	VSS	4.00835e-17	$cmodel
C23	BL<28>	VSS	4.00324e-17	$cmodel
C24	BL<29>	VSS	4.00835e-17	$cmodel
C25	BL<2>	VSS	4.00324e-17	$cmodel
C26	BL<30>	VSS	4.00324e-17	$cmodel
C27	BL<31>	VSS	4.00835e-17	$cmodel
C28	BL<32>	VSS	4.00324e-17	$cmodel
C29	BL<33>	VSS	4.00835e-17	$cmodel
C30	BL<34>	VSS	4.00324e-17	$cmodel
C31	BL<35>	VSS	4.00835e-17	$cmodel
C32	BL<36>	VSS	4.00324e-17	$cmodel
C33	BL<37>	VSS	4.00835e-17	$cmodel
C34	BL<38>	VSS	4.00324e-17	$cmodel
C35	BL<39>	VSS	4.00835e-17	$cmodel
C36	BL<3>	VSS	4.00835e-17	$cmodel
C37	BL<40>	VSS	4.00324e-17	$cmodel
C38	BL<41>	VSS	4.00835e-17	$cmodel
C39	BL<42>	VSS	4.00324e-17	$cmodel
C40	BL<43>	VSS	4.00835e-17	$cmodel
C41	BL<44>	VSS	4.00324e-17	$cmodel
C42	BL<45>	VSS	4.00835e-17	$cmodel
C43	BL<46>	VSS	4.00324e-17	$cmodel
C44	BL<47>	VSS	4.00835e-17	$cmodel
C45	BL<48>	VSS	4.00324e-17	$cmodel
C46	BL<49>	VSS	4.00835e-17	$cmodel
C47	BL<4>	VSS	4.00324e-17	$cmodel
C48	BL<50>	VSS	4.00324e-17	$cmodel
C49	BL<51>	VSS	4.00835e-17	$cmodel
C50	BL<52>	VSS	4.00324e-17	$cmodel
C51	BL<53>	VSS	4.00835e-17	$cmodel
C52	BL<54>	VSS	4.00324e-17	$cmodel
C53	BL<55>	VSS	4.00835e-17	$cmodel
C54	BL<56>	VSS	4.00324e-17	$cmodel
C55	BL<57>	VSS	4.00835e-17	$cmodel
C56	BL<58>	VSS	4.00324e-17	$cmodel
C57	BL<59>	VSS	4.00835e-17	$cmodel
C58	BL<5>	VSS	4.00835e-17	$cmodel
C59	BL<60>	VSS	4.00324e-17	$cmodel
C60	BL<61>	VSS	4.00835e-17	$cmodel
C61	BL<62>	VSS	4.00324e-17	$cmodel
C62	BL<63>	VSS	4.1541e-17	$cmodel
C63	BL<6>	VSS	4.00324e-17	$cmodel
C64	BL<7>	VSS	4.00835e-17	$cmodel
C65	BL<8>	VSS	4.00324e-17	$cmodel
C66	BL<9>	VSS	4.00835e-17	$cmodel
C67	BLB<0>	VSS	1.4668e-17	$cmodel
C68	BLB<10>	VSS	1.4668e-17	$cmodel
C69	BLB<11>	VSS	1.4668e-17	$cmodel
C70	BLB<12>	VSS	1.4668e-17	$cmodel
C71	BLB<13>	VSS	1.4668e-17	$cmodel
C72	BLB<14>	VSS	1.4668e-17	$cmodel
C73	BLB<15>	VSS	1.4668e-17	$cmodel
C74	BLB<16>	VSS	1.4668e-17	$cmodel
C75	BLB<17>	VSS	1.4668e-17	$cmodel
C76	BLB<18>	VSS	1.4668e-17	$cmodel
C77	BLB<19>	VSS	1.4668e-17	$cmodel
C78	BLB<1>	VSS	1.4668e-17	$cmodel
C79	BLB<20>	VSS	1.4668e-17	$cmodel
C80	BLB<21>	VSS	1.4668e-17	$cmodel
C81	BLB<22>	VSS	1.4668e-17	$cmodel
C82	BLB<23>	VSS	1.4668e-17	$cmodel
C83	BLB<24>	VSS	1.4668e-17	$cmodel
C84	BLB<25>	VSS	1.4668e-17	$cmodel
C85	BLB<26>	VSS	1.4668e-17	$cmodel
C86	BLB<27>	VSS	1.4668e-17	$cmodel
C87	BLB<28>	VSS	1.4668e-17	$cmodel
C88	BLB<29>	VSS	1.4668e-17	$cmodel
C89	BLB<2>	VSS	1.4668e-17	$cmodel
C90	BLB<30>	VSS	1.4668e-17	$cmodel
C91	BLB<31>	VSS	1.4668e-17	$cmodel
C92	BLB<32>	VSS	1.4668e-17	$cmodel
C93	BLB<33>	VSS	1.4668e-17	$cmodel
C94	BLB<34>	VSS	1.4668e-17	$cmodel
C95	BLB<35>	VSS	1.4668e-17	$cmodel
C96	BLB<36>	VSS	1.4668e-17	$cmodel
C97	BLB<37>	VSS	1.4668e-17	$cmodel
C98	BLB<38>	VSS	1.4668e-17	$cmodel
C99	BLB<39>	VSS	1.4668e-17	$cmodel
C100	BLB<3>	VSS	1.4668e-17	$cmodel
C101	BLB<40>	VSS	1.4668e-17	$cmodel
C102	BLB<41>	VSS	1.4668e-17	$cmodel
C103	BLB<42>	VSS	1.4668e-17	$cmodel
C104	BLB<43>	VSS	1.4668e-17	$cmodel
C105	BLB<44>	VSS	1.4668e-17	$cmodel
C106	BLB<45>	VSS	1.4668e-17	$cmodel
C107	BLB<46>	VSS	1.4668e-17	$cmodel
C108	BLB<47>	VSS	1.4668e-17	$cmodel
C109	BLB<48>	VSS	1.4668e-17	$cmodel
C110	BLB<49>	VSS	1.4668e-17	$cmodel
C111	BLB<4>	VSS	1.4668e-17	$cmodel
C112	BLB<50>	VSS	1.4668e-17	$cmodel
C113	BLB<51>	VSS	1.4668e-17	$cmodel
C114	BLB<52>	VSS	1.4668e-17	$cmodel
C115	BLB<53>	VSS	1.4668e-17	$cmodel
C116	BLB<54>	VSS	1.4668e-17	$cmodel
C117	BLB<55>	VSS	1.4668e-17	$cmodel
C118	BLB<56>	VSS	1.4668e-17	$cmodel
C119	BLB<57>	VSS	1.4668e-17	$cmodel
C120	BLB<58>	VSS	1.4668e-17	$cmodel
C121	BLB<59>	VSS	1.4668e-17	$cmodel
C122	BLB<5>	VSS	1.4668e-17	$cmodel
C123	BLB<60>	VSS	1.4668e-17	$cmodel
C124	BLB<61>	VSS	1.4668e-17	$cmodel
C125	BLB<62>	VSS	1.4668e-17	$cmodel
C126	BLB<63>	VSS	1.61489e-17	$cmodel
C127	BLB<6>	VSS	1.4668e-17	$cmodel
C128	BLB<7>	VSS	1.4668e-17	$cmodel
C129	BLB<8>	VSS	1.4668e-17	$cmodel
C130	BLB<9>	VSS	1.4668e-17	$cmodel
C131	I0<7>/I1<7>/QB	VSS	4.18748e-17	$cmodel
C132	I0<7>/I1<7>/Q	VSS	7.79049e-17	$cmodel
C133	I0<7>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C134	I0<7>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C135	I0<7>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C136	I0<7>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C137	I0<7>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C138	I0<7>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C139	I0<7>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C140	I0<7>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C141	I0<7>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C142	I0<7>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C143	I0<7>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C144	I0<7>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C145	I0<7>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C146	I0<7>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C147	I0<6>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C148	I0<6>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C149	I0<6>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C150	I0<6>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C151	I0<6>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C152	I0<6>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C153	I0<6>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C154	I0<6>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C155	I0<6>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C156	I0<6>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C157	I0<6>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C158	I0<6>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C159	I0<6>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C160	I0<6>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C161	I0<6>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C162	I0<6>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C163	I0<5>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C164	I0<5>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C165	I0<5>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C166	I0<5>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C167	I0<5>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C168	I0<5>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C169	I0<5>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C170	I0<5>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C171	I0<5>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C172	I0<5>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C173	I0<5>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C174	I0<5>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C175	I0<5>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C176	I0<5>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C177	I0<5>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C178	I0<5>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C179	I0<4>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C180	I0<4>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C181	I0<4>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C182	I0<4>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C183	I0<4>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C184	I0<4>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C185	I0<4>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C186	I0<4>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C187	I0<4>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C188	I0<4>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C189	I0<4>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C190	I0<4>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C191	I0<4>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C192	I0<4>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C193	I0<4>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C194	I0<4>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C195	I0<3>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C196	I0<3>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C197	I0<3>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C198	I0<3>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C199	I0<3>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C200	I0<3>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C201	I0<3>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C202	I0<3>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C203	I0<3>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C204	I0<3>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C205	I0<3>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C206	I0<3>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C207	I0<3>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C208	I0<3>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C209	I0<3>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C210	I0<3>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C211	I0<2>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C212	I0<2>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C213	I0<2>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C214	I0<2>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C215	I0<2>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C216	I0<2>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C217	I0<2>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C218	I0<2>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C219	I0<2>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C220	I0<2>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C221	I0<2>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C222	I0<2>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C223	I0<2>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C224	I0<2>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C225	I0<2>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C226	I0<2>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C227	I0<1>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C228	I0<1>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C229	I0<1>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C230	I0<1>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C231	I0<1>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C232	I0<1>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C233	I0<1>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C234	I0<1>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C235	I0<1>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C236	I0<1>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C237	I0<1>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C238	I0<1>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C239	I0<1>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C240	I0<1>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C241	I0<1>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C242	I0<1>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C243	I0<0>/I1<7>/QB	VSS	3.96263e-17	$cmodel
C244	I0<0>/I1<7>/Q	VSS	7.7884e-17	$cmodel
C245	I0<0>/I1<6>/QB	VSS	3.96263e-17	$cmodel
C246	I0<0>/I1<6>/Q	VSS	7.7884e-17	$cmodel
C247	I0<0>/I1<5>/QB	VSS	2.18331e-17	$cmodel
C248	I0<0>/I1<5>/Q	VSS	4.19596e-17	$cmodel
C249	I0<0>/I1<4>/QB	VSS	3.96263e-17	$cmodel
C250	I0<0>/I1<4>/Q	VSS	7.7884e-17	$cmodel
C251	I0<0>/I1<3>/QB	VSS	2.18331e-17	$cmodel
C252	I0<0>/I1<3>/Q	VSS	4.19596e-17	$cmodel
C253	I0<0>/I1<2>/QB	VSS	3.96263e-17	$cmodel
C254	I0<0>/I1<2>/Q	VSS	7.7884e-17	$cmodel
C255	I0<0>/I1<1>/QB	VSS	2.18331e-17	$cmodel
C256	I0<0>/I1<1>/Q	VSS	4.19596e-17	$cmodel
C257	I0<0>/I1<0>/QB	VSS	2.18331e-17	$cmodel
C258	I0<0>/I1<0>/Q	VSS	4.19596e-17	$cmodel
C259	I0<7>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C260	I0<7>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C261	I0<7>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C262	I0<7>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C263	I0<7>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C264	I0<7>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C265	I0<7>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C266	I0<7>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C267	I0<7>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C268	I0<7>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C269	I0<7>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C270	I0<7>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C271	I0<6>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C272	I0<6>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C273	I0<6>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C274	I0<6>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C275	I0<6>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C276	I0<6>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C277	I0<6>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C278	I0<6>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C279	I0<6>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C280	I0<6>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C281	I0<6>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C282	I0<6>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C283	I0<5>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C284	I0<5>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C285	I0<5>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C286	I0<5>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C287	I0<5>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C288	I0<5>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C289	I0<5>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C290	I0<5>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C291	I0<5>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C292	I0<5>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C293	I0<5>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C294	I0<5>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C295	I0<4>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C296	I0<4>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C297	I0<4>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C298	I0<4>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C299	I0<4>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C300	I0<4>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C301	I0<4>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C302	I0<4>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C303	I0<4>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C304	I0<4>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C305	I0<4>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C306	I0<4>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C307	I0<3>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C308	I0<3>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C309	I0<3>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C310	I0<3>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C311	I0<3>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C312	I0<3>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C313	I0<3>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C314	I0<3>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C315	I0<3>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C316	I0<3>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C317	I0<3>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C318	I0<3>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C319	I0<2>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C320	I0<2>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C321	I0<2>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C322	I0<2>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C323	I0<2>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C324	I0<2>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C325	I0<2>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C326	I0<2>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C327	I0<2>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C328	I0<2>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C329	I0<2>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C330	I0<2>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C331	I0<1>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C332	I0<1>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C333	I0<1>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C334	I0<1>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C335	I0<1>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C336	I0<1>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C337	I0<1>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C338	I0<1>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C339	I0<1>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C340	I0<1>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C341	I0<1>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C342	I0<1>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C343	I0<0>/I1<7>/QB#2	VSS	2.19709e-17	$cmodel
C344	I0<0>/I1<7>/Q#2	VSS	2.421e-17	$cmodel
C345	I0<0>/I1<5>/Q#2	VSS	2.4257e-17	$cmodel
C346	I0<0>/I1<6>/QB#2	VSS	2.19709e-17	$cmodel
C347	I0<0>/I1<6>/Q#2	VSS	2.421e-17	$cmodel
C348	I0<0>/I1<3>/Q#2	VSS	2.4257e-17	$cmodel
C349	I0<0>/I1<4>/QB#2	VSS	2.19709e-17	$cmodel
C350	I0<0>/I1<4>/Q#2	VSS	2.421e-17	$cmodel
C351	I0<0>/I1<1>/Q#2	VSS	2.4257e-17	$cmodel
C352	I0<0>/I1<2>/QB#2	VSS	2.19709e-17	$cmodel
C353	I0<0>/I1<2>/Q#2	VSS	2.421e-17	$cmodel
C354	I0<0>/I1<0>/Q#2	VSS	2.4257e-17	$cmodel
C355	WL#254	VSS	2.94557e-17	$cmodel
C356	I0<7>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C357	WL#250	VSS	2.91904e-17	$cmodel
C358	WL#252	VSS	2.89999e-17	$cmodel
C359	WL#246	VSS	2.96063e-17	$cmodel
C360	I0<7>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C361	WL#248	VSS	2.95464e-17	$cmodel
C362	I0<7>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C363	WL#242	VSS	2.91904e-17	$cmodel
C364	WL#244	VSS	2.89999e-17	$cmodel
C365	WL#238	VSS	2.96063e-17	$cmodel
C366	I0<7>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C367	WL#240	VSS	2.95464e-17	$cmodel
C368	I0<7>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C369	WL#234	VSS	2.91904e-17	$cmodel
C370	WL#236	VSS	2.89999e-17	$cmodel
C371	WL#230	VSS	2.96063e-17	$cmodel
C372	I0<7>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C373	WL#232	VSS	2.95464e-17	$cmodel
C374	I0<7>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C375	WL#226	VSS	2.91904e-17	$cmodel
C376	WL#228	VSS	2.89999e-17	$cmodel
C377	WL#222	VSS	2.96063e-17	$cmodel
C378	I0<7>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C379	WL#224	VSS	2.95464e-17	$cmodel
C380	I0<6>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C381	WL#218	VSS	2.91904e-17	$cmodel
C382	WL#220	VSS	2.89999e-17	$cmodel
C383	WL#214	VSS	2.96063e-17	$cmodel
C384	I0<6>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C385	WL#216	VSS	2.95464e-17	$cmodel
C386	I0<6>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C387	WL#210	VSS	2.91904e-17	$cmodel
C388	WL#212	VSS	2.89999e-17	$cmodel
C389	WL#206	VSS	2.96063e-17	$cmodel
C390	I0<6>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C391	WL#208	VSS	2.95464e-17	$cmodel
C392	I0<6>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C393	WL#202	VSS	2.91904e-17	$cmodel
C394	WL#204	VSS	2.89999e-17	$cmodel
C395	WL#198	VSS	2.96063e-17	$cmodel
C396	I0<6>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C397	WL#200	VSS	2.95464e-17	$cmodel
C398	I0<6>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C399	WL#194	VSS	2.91904e-17	$cmodel
C400	WL#196	VSS	2.89999e-17	$cmodel
C401	WL#190	VSS	2.96063e-17	$cmodel
C402	I0<6>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C403	WL#192	VSS	2.95464e-17	$cmodel
C404	I0<5>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C405	WL#186	VSS	2.91904e-17	$cmodel
C406	WL#188	VSS	2.89999e-17	$cmodel
C407	WL#182	VSS	2.96063e-17	$cmodel
C408	I0<5>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C409	WL#184	VSS	2.95464e-17	$cmodel
C410	I0<5>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C411	WL#178	VSS	2.91904e-17	$cmodel
C412	WL#180	VSS	2.89999e-17	$cmodel
C413	WL#174	VSS	2.96063e-17	$cmodel
C414	I0<5>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C415	WL#176	VSS	2.95464e-17	$cmodel
C416	I0<5>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C417	WL#170	VSS	2.91904e-17	$cmodel
C418	WL#172	VSS	2.89999e-17	$cmodel
C419	WL#166	VSS	2.96063e-17	$cmodel
C420	I0<5>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C421	WL#168	VSS	2.95464e-17	$cmodel
C422	I0<5>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C423	WL#162	VSS	2.91904e-17	$cmodel
C424	WL#164	VSS	2.89999e-17	$cmodel
C425	WL#158	VSS	2.96063e-17	$cmodel
C426	I0<5>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C427	WL#160	VSS	2.95464e-17	$cmodel
C428	I0<4>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C429	WL#154	VSS	2.91904e-17	$cmodel
C430	WL#156	VSS	2.89999e-17	$cmodel
C431	WL#150	VSS	2.96063e-17	$cmodel
C432	I0<4>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C433	WL#152	VSS	2.95464e-17	$cmodel
C434	I0<4>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C435	WL#146	VSS	2.91904e-17	$cmodel
C436	WL#148	VSS	2.89999e-17	$cmodel
C437	WL#142	VSS	2.96063e-17	$cmodel
C438	I0<4>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C439	WL#144	VSS	2.95464e-17	$cmodel
C440	I0<4>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C441	WL#138	VSS	2.91904e-17	$cmodel
C442	WL#140	VSS	2.89999e-17	$cmodel
C443	WL#134	VSS	2.96063e-17	$cmodel
C444	I0<4>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C445	WL#136	VSS	2.95464e-17	$cmodel
C446	I0<4>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C447	WL#130	VSS	2.91904e-17	$cmodel
C448	WL#132	VSS	2.89999e-17	$cmodel
C449	WL#126	VSS	2.96063e-17	$cmodel
C450	I0<4>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C451	WL#128	VSS	2.95464e-17	$cmodel
C452	I0<3>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C453	WL#122	VSS	2.91904e-17	$cmodel
C454	WL#124	VSS	2.89999e-17	$cmodel
C455	WL#118	VSS	2.96063e-17	$cmodel
C456	I0<3>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C457	WL#120	VSS	2.95464e-17	$cmodel
C458	I0<3>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C459	WL#114	VSS	2.91904e-17	$cmodel
C460	WL#116	VSS	2.89999e-17	$cmodel
C461	WL#110	VSS	2.96063e-17	$cmodel
C462	I0<3>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C463	WL#112	VSS	2.95464e-17	$cmodel
C464	I0<3>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C465	WL#106	VSS	2.91904e-17	$cmodel
C466	WL#108	VSS	2.89999e-17	$cmodel
C467	WL#102	VSS	2.96063e-17	$cmodel
C468	I0<3>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C469	WL#104	VSS	2.95464e-17	$cmodel
C470	I0<3>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C471	WL#98	VSS	2.91904e-17	$cmodel
C472	WL#100	VSS	2.89999e-17	$cmodel
C473	WL#94	VSS	2.96063e-17	$cmodel
C474	I0<3>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C475	WL#96	VSS	2.95464e-17	$cmodel
C476	I0<2>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C477	WL#90	VSS	2.91904e-17	$cmodel
C478	WL#92	VSS	2.89999e-17	$cmodel
C479	WL#86	VSS	2.96063e-17	$cmodel
C480	I0<2>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C481	WL#88	VSS	2.95464e-17	$cmodel
C482	I0<2>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C483	WL#82	VSS	2.91904e-17	$cmodel
C484	WL#84	VSS	2.89999e-17	$cmodel
C485	WL#78	VSS	2.96063e-17	$cmodel
C486	I0<2>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C487	WL#80	VSS	2.95464e-17	$cmodel
C488	I0<2>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C489	WL#74	VSS	2.91904e-17	$cmodel
C490	WL#76	VSS	2.89999e-17	$cmodel
C491	WL#70	VSS	2.96063e-17	$cmodel
C492	I0<2>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C493	WL#72	VSS	2.95464e-17	$cmodel
C494	I0<2>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C495	WL#66	VSS	2.91904e-17	$cmodel
C496	WL#68	VSS	2.89999e-17	$cmodel
C497	WL#62	VSS	2.96063e-17	$cmodel
C498	I0<2>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C499	WL#64	VSS	2.95464e-17	$cmodel
C500	I0<1>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C501	WL#58	VSS	2.91904e-17	$cmodel
C502	WL#60	VSS	2.89999e-17	$cmodel
C503	WL#54	VSS	2.96063e-17	$cmodel
C504	I0<1>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C505	WL#56	VSS	2.95464e-17	$cmodel
C506	I0<1>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C507	WL#50	VSS	2.91904e-17	$cmodel
C508	WL#52	VSS	2.89999e-17	$cmodel
C509	WL#46	VSS	2.96063e-17	$cmodel
C510	I0<1>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C511	WL#48	VSS	2.95464e-17	$cmodel
C512	I0<1>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C513	WL#42	VSS	2.91904e-17	$cmodel
C514	WL#44	VSS	2.89999e-17	$cmodel
C515	WL#38	VSS	2.96063e-17	$cmodel
C516	I0<1>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C517	WL#40	VSS	2.95464e-17	$cmodel
C518	I0<1>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C519	WL#34	VSS	2.91904e-17	$cmodel
C520	WL#36	VSS	2.89999e-17	$cmodel
C521	WL#30	VSS	2.96063e-17	$cmodel
C522	I0<1>/I1<0>/QB#2	VSS	3.97013e-17	$cmodel
C523	WL#32	VSS	2.95464e-17	$cmodel
C524	I0<0>/I1<7>/Q#3	VSS	4.24109e-17	$cmodel
C525	WL#26	VSS	2.91904e-17	$cmodel
C526	WL#28	VSS	2.89999e-17	$cmodel
C527	WL#22	VSS	2.96063e-17	$cmodel
C528	I0<0>/I1<5>/QB#2	VSS	3.97013e-17	$cmodel
C529	WL#24	VSS	2.95464e-17	$cmodel
C530	I0<0>/I1<6>/Q#3	VSS	4.24109e-17	$cmodel
C531	WL#18	VSS	2.91904e-17	$cmodel
C532	WL#20	VSS	2.89999e-17	$cmodel
C533	WL#14	VSS	2.96063e-17	$cmodel
C534	I0<0>/I1<3>/QB#2	VSS	3.97013e-17	$cmodel
C535	WL#16	VSS	2.95464e-17	$cmodel
C536	I0<0>/I1<4>/Q#3	VSS	4.24109e-17	$cmodel
C537	WL#10	VSS	2.91904e-17	$cmodel
C538	WL#12	VSS	2.89999e-17	$cmodel
C539	WL#6	VSS	2.96063e-17	$cmodel
C540	I0<0>/I1<1>/QB#2	VSS	3.97013e-17	$cmodel
C541	WL#8	VSS	2.95464e-17	$cmodel
C542	I0<0>/I1<2>/Q#3	VSS	4.24109e-17	$cmodel
C543	WL#3	VSS	2.91904e-17	$cmodel
C544	WL#5	VSS	2.89999e-17	$cmodel
C545	WL#1	VSS	2.95243e-17	$cmodel
C546	I0<0>/I1<0>/QB#2	VSS	4.19392e-17	$cmodel
C547	WL#255	VSS	2.94109e-17	$cmodel
C548	I0<7>/I1<7>/QB#3	VSS	7.92335e-17	$cmodel
C549	WL#251	VSS	3.01301e-17	$cmodel
C550	I0<7>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C551	I0<7>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C552	WL#247	VSS	3.68326e-17	$cmodel
C553	I0<7>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C554	WL#243	VSS	3.01464e-17	$cmodel
C555	I0<7>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C556	I0<7>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C557	WL#239	VSS	3.68326e-17	$cmodel
C558	I0<7>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C559	WL#235	VSS	3.01464e-17	$cmodel
C560	I0<7>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C561	I0<7>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C562	WL#231	VSS	3.68326e-17	$cmodel
C563	I0<7>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C564	WL#227	VSS	3.01464e-17	$cmodel
C565	I0<7>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C566	I0<7>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C567	WL#223	VSS	3.68326e-17	$cmodel
C568	I0<6>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C569	WL#219	VSS	3.01464e-17	$cmodel
C570	I0<6>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C571	I0<6>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C572	WL#215	VSS	3.68326e-17	$cmodel
C573	I0<6>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C574	WL#211	VSS	3.01464e-17	$cmodel
C575	I0<6>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C576	I0<6>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C577	WL#207	VSS	3.68326e-17	$cmodel
C578	I0<6>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C579	WL#203	VSS	3.01464e-17	$cmodel
C580	I0<6>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C581	I0<6>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C582	WL#199	VSS	3.68326e-17	$cmodel
C583	I0<6>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C584	WL#195	VSS	3.01464e-17	$cmodel
C585	I0<6>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C586	I0<6>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C587	WL#191	VSS	3.68326e-17	$cmodel
C588	I0<5>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C589	WL#187	VSS	3.01464e-17	$cmodel
C590	I0<5>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C591	I0<5>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C592	WL#183	VSS	3.68326e-17	$cmodel
C593	I0<5>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C594	WL#179	VSS	3.01464e-17	$cmodel
C595	I0<5>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C596	I0<5>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C597	WL#175	VSS	3.68326e-17	$cmodel
C598	I0<5>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C599	WL#171	VSS	3.01464e-17	$cmodel
C600	I0<5>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C601	I0<5>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C602	WL#167	VSS	3.68326e-17	$cmodel
C603	I0<5>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C604	WL#163	VSS	3.01464e-17	$cmodel
C605	I0<5>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C606	I0<5>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C607	WL#159	VSS	3.68326e-17	$cmodel
C608	I0<4>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C609	WL#155	VSS	3.01464e-17	$cmodel
C610	I0<4>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C611	I0<4>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C612	WL#151	VSS	3.68326e-17	$cmodel
C613	I0<4>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C614	WL#147	VSS	3.01464e-17	$cmodel
C615	I0<4>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C616	I0<4>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C617	WL#143	VSS	3.68326e-17	$cmodel
C618	I0<4>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C619	WL#139	VSS	3.01464e-17	$cmodel
C620	I0<4>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C621	I0<4>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C622	WL#135	VSS	3.68326e-17	$cmodel
C623	I0<4>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C624	WL#131	VSS	3.01464e-17	$cmodel
C625	I0<4>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C626	I0<4>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C627	WL#127	VSS	3.68326e-17	$cmodel
C628	I0<3>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C629	WL#123	VSS	3.01464e-17	$cmodel
C630	I0<3>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C631	I0<3>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C632	WL#119	VSS	3.68326e-17	$cmodel
C633	I0<3>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C634	WL#115	VSS	3.01464e-17	$cmodel
C635	I0<3>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C636	I0<3>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C637	WL#111	VSS	3.68326e-17	$cmodel
C638	I0<3>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C639	WL#107	VSS	3.01464e-17	$cmodel
C640	I0<3>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C641	I0<3>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C642	WL#103	VSS	3.68326e-17	$cmodel
C643	I0<3>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C644	WL#99	VSS	3.01464e-17	$cmodel
C645	I0<3>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C646	I0<3>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C647	WL#95	VSS	3.68326e-17	$cmodel
C648	I0<2>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C649	WL#91	VSS	3.01464e-17	$cmodel
C650	I0<2>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C651	I0<2>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C652	WL#87	VSS	3.68326e-17	$cmodel
C653	I0<2>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C654	WL#83	VSS	3.01464e-17	$cmodel
C655	I0<2>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C656	I0<2>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C657	WL#79	VSS	3.68326e-17	$cmodel
C658	I0<2>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C659	WL#75	VSS	3.01464e-17	$cmodel
C660	I0<2>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C661	I0<2>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C662	WL#71	VSS	3.68326e-17	$cmodel
C663	I0<2>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C664	WL#67	VSS	3.01464e-17	$cmodel
C665	I0<2>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C666	I0<2>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C667	WL#63	VSS	3.68326e-17	$cmodel
C668	I0<1>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C669	WL#59	VSS	3.01464e-17	$cmodel
C670	I0<1>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C671	I0<1>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C672	WL#55	VSS	3.68326e-17	$cmodel
C673	I0<1>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C674	WL#51	VSS	3.01464e-17	$cmodel
C675	I0<1>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C676	I0<1>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C677	WL#47	VSS	3.68326e-17	$cmodel
C678	I0<1>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C679	WL#43	VSS	3.01464e-17	$cmodel
C680	I0<1>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C681	I0<1>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C682	WL#39	VSS	3.68326e-17	$cmodel
C683	I0<1>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C684	WL#35	VSS	3.01464e-17	$cmodel
C685	I0<1>/I1<0>/QB#3	VSS	8.01335e-17	$cmodel
C686	I0<1>/I1<0>/Q#3	VSS	7.64904e-17	$cmodel
C687	WL#31	VSS	3.68326e-17	$cmodel
C688	I0<0>/I1<7>/QB#3	VSS	7.94925e-17	$cmodel
C689	WL#27	VSS	3.01464e-17	$cmodel
C690	I0<0>/I1<5>/QB#3	VSS	8.01335e-17	$cmodel
C691	I0<0>/I1<5>/Q#3	VSS	7.64904e-17	$cmodel
C692	WL#23	VSS	3.68326e-17	$cmodel
C693	I0<0>/I1<6>/QB#3	VSS	7.94925e-17	$cmodel
C694	WL#19	VSS	3.01464e-17	$cmodel
C695	I0<0>/I1<3>/QB#3	VSS	8.01335e-17	$cmodel
C696	I0<0>/I1<3>/Q#3	VSS	7.64904e-17	$cmodel
C697	WL#15	VSS	3.68326e-17	$cmodel
C698	I0<0>/I1<4>/QB#3	VSS	7.94925e-17	$cmodel
C699	WL#11	VSS	3.01464e-17	$cmodel
C700	I0<0>/I1<1>/QB#3	VSS	8.01335e-17	$cmodel
C701	I0<0>/I1<1>/Q#3	VSS	7.64904e-17	$cmodel
C702	WL#7	VSS	3.68326e-17	$cmodel
C703	I0<0>/I1<2>/QB#3	VSS	7.94925e-17	$cmodel
C704	WL#4	VSS	3.01423e-17	$cmodel
C705	I0<0>/I1<0>/QB#3	VSS	7.9902e-17	$cmodel
C706	I0<0>/I1<0>/Q#3	VSS	7.65082e-17	$cmodel
C707	WL#2	VSS	2.7968e-17	$cmodel
C708	BL<63>#3	VSS	8.79767e-17	$cmodel
C709	VDD#572	VSS	2.50983e-17	$cmodel
C710	VDD#573	VSS	2.04193e-17	$cmodel
C711	BLB<63>#3	VSS	1.28005e-16	$cmodel
C712	BLB<62>#3	VSS	7.41005e-17	$cmodel
C713	VDD#570	VSS	5.91314e-17	$cmodel
C714	VDD#571	VSS	5.94258e-17	$cmodel
C715	BL<62>#3	VSS	4.79226e-17	$cmodel
C716	BL<61>#3	VSS	8.82729e-17	$cmodel
C717	VDD#568	VSS	2.49053e-17	$cmodel
C718	VDD#569	VSS	2.50001e-17	$cmodel
C719	BLB<61>#3	VSS	1.28016e-16	$cmodel
C720	BLB<60>#2	VSS	7.41074e-17	$cmodel
C721	VDD#547	VSS	5.91314e-17	$cmodel
C722	VDD#548	VSS	5.94258e-17	$cmodel
C723	BL<60>#3	VSS	4.79226e-17	$cmodel
C724	BL<59>#3	VSS	8.82729e-17	$cmodel
C725	VDD#538	VSS	2.49053e-17	$cmodel
C726	VDD#539	VSS	2.50001e-17	$cmodel
C727	BLB<59>#3	VSS	1.28016e-16	$cmodel
C728	BLB<58>#2	VSS	7.41074e-17	$cmodel
C729	VDD#529	VSS	5.91314e-17	$cmodel
C730	VDD#530	VSS	5.94258e-17	$cmodel
C731	BL<58>#3	VSS	4.79226e-17	$cmodel
C732	BL<57>#3	VSS	8.82729e-17	$cmodel
C733	VDD#520	VSS	2.49053e-17	$cmodel
C734	VDD#521	VSS	2.50001e-17	$cmodel
C735	BLB<57>#3	VSS	1.28016e-16	$cmodel
C736	BLB<56>#2	VSS	7.41074e-17	$cmodel
C737	VDD#511	VSS	5.91314e-17	$cmodel
C738	VDD#512	VSS	5.94258e-17	$cmodel
C739	BL<56>#3	VSS	4.79226e-17	$cmodel
C740	BL<55>#3	VSS	8.82729e-17	$cmodel
C741	VDD#502	VSS	2.49053e-17	$cmodel
C742	VDD#503	VSS	2.50001e-17	$cmodel
C743	BLB<55>#3	VSS	1.28016e-16	$cmodel
C744	BLB<54>#2	VSS	7.41074e-17	$cmodel
C745	VDD#493	VSS	5.91314e-17	$cmodel
C746	VDD#494	VSS	5.94258e-17	$cmodel
C747	BL<54>#3	VSS	4.79226e-17	$cmodel
C748	BL<53>#3	VSS	8.82729e-17	$cmodel
C749	VDD#484	VSS	2.49053e-17	$cmodel
C750	VDD#485	VSS	2.50001e-17	$cmodel
C751	BLB<53>#3	VSS	1.28016e-16	$cmodel
C752	BLB<52>#2	VSS	7.41074e-17	$cmodel
C753	VDD#475	VSS	5.91314e-17	$cmodel
C754	VDD#476	VSS	5.94258e-17	$cmodel
C755	BL<52>#3	VSS	4.79226e-17	$cmodel
C756	BL<51>#3	VSS	8.82729e-17	$cmodel
C757	VDD#466	VSS	2.49053e-17	$cmodel
C758	VDD#467	VSS	2.50001e-17	$cmodel
C759	BLB<51>#3	VSS	1.28016e-16	$cmodel
C760	BLB<50>#2	VSS	7.41074e-17	$cmodel
C761	VDD#457	VSS	5.91314e-17	$cmodel
C762	VDD#458	VSS	5.94258e-17	$cmodel
C763	BL<50>#3	VSS	4.79226e-17	$cmodel
C764	BL<49>#3	VSS	8.82729e-17	$cmodel
C765	VDD#448	VSS	2.49053e-17	$cmodel
C766	VDD#449	VSS	2.50001e-17	$cmodel
C767	BLB<49>#3	VSS	1.28016e-16	$cmodel
C768	BLB<48>#2	VSS	7.41074e-17	$cmodel
C769	VDD#439	VSS	5.91314e-17	$cmodel
C770	VDD#440	VSS	5.94258e-17	$cmodel
C771	BL<48>#3	VSS	4.79226e-17	$cmodel
C772	BL<47>#3	VSS	8.82729e-17	$cmodel
C773	VDD#430	VSS	2.49053e-17	$cmodel
C774	VDD#431	VSS	2.50001e-17	$cmodel
C775	BLB<47>#3	VSS	1.28016e-16	$cmodel
C776	BLB<46>#2	VSS	7.41074e-17	$cmodel
C777	VDD#421	VSS	5.91314e-17	$cmodel
C778	VDD#422	VSS	5.94258e-17	$cmodel
C779	BL<46>#3	VSS	4.79226e-17	$cmodel
C780	BL<45>#3	VSS	8.82729e-17	$cmodel
C781	VDD#412	VSS	2.49053e-17	$cmodel
C782	VDD#413	VSS	2.50001e-17	$cmodel
C783	BLB<45>#3	VSS	1.28016e-16	$cmodel
C784	BLB<44>#2	VSS	7.41074e-17	$cmodel
C785	VDD#403	VSS	5.91314e-17	$cmodel
C786	VDD#404	VSS	5.94258e-17	$cmodel
C787	BL<44>#3	VSS	4.79226e-17	$cmodel
C788	BL<43>#3	VSS	8.82729e-17	$cmodel
C789	VDD#394	VSS	2.49053e-17	$cmodel
C790	VDD#395	VSS	2.50001e-17	$cmodel
C791	BLB<43>#3	VSS	1.28016e-16	$cmodel
C792	BLB<42>#2	VSS	7.41074e-17	$cmodel
C793	VDD#385	VSS	5.91314e-17	$cmodel
C794	VDD#386	VSS	5.94258e-17	$cmodel
C795	BL<42>#3	VSS	4.79226e-17	$cmodel
C796	BL<41>#3	VSS	8.82729e-17	$cmodel
C797	VDD#376	VSS	2.49053e-17	$cmodel
C798	VDD#377	VSS	2.50001e-17	$cmodel
C799	BLB<41>#3	VSS	1.28016e-16	$cmodel
C800	BLB<40>#2	VSS	7.41074e-17	$cmodel
C801	VDD#367	VSS	5.91314e-17	$cmodel
C802	VDD#368	VSS	5.94258e-17	$cmodel
C803	BL<40>#3	VSS	4.79226e-17	$cmodel
C804	BL<39>#3	VSS	8.82729e-17	$cmodel
C805	VDD#358	VSS	2.49053e-17	$cmodel
C806	VDD#359	VSS	2.50001e-17	$cmodel
C807	BLB<39>#3	VSS	1.28016e-16	$cmodel
C808	BLB<38>#2	VSS	7.41074e-17	$cmodel
C809	VDD#349	VSS	5.91314e-17	$cmodel
C810	VDD#350	VSS	5.94258e-17	$cmodel
C811	BL<38>#3	VSS	4.79226e-17	$cmodel
C812	BL<37>#3	VSS	8.82729e-17	$cmodel
C813	VDD#340	VSS	2.49053e-17	$cmodel
C814	VDD#341	VSS	2.50001e-17	$cmodel
C815	BLB<37>#3	VSS	1.28016e-16	$cmodel
C816	BLB<36>#2	VSS	7.41074e-17	$cmodel
C817	VDD#331	VSS	5.91314e-17	$cmodel
C818	VDD#332	VSS	5.94258e-17	$cmodel
C819	BL<36>#3	VSS	4.79226e-17	$cmodel
C820	BL<35>#3	VSS	8.82729e-17	$cmodel
C821	VDD#322	VSS	2.49053e-17	$cmodel
C822	VDD#323	VSS	2.50001e-17	$cmodel
C823	BLB<35>#3	VSS	1.28016e-16	$cmodel
C824	BLB<34>#2	VSS	7.41074e-17	$cmodel
C825	VDD#313	VSS	5.91314e-17	$cmodel
C826	VDD#314	VSS	5.94258e-17	$cmodel
C827	BL<34>#3	VSS	4.79226e-17	$cmodel
C828	BL<33>#3	VSS	8.82729e-17	$cmodel
C829	VDD#304	VSS	2.49053e-17	$cmodel
C830	VDD#305	VSS	2.50001e-17	$cmodel
C831	BLB<33>#3	VSS	1.28016e-16	$cmodel
C832	BLB<32>#2	VSS	7.41074e-17	$cmodel
C833	VDD#295	VSS	5.91314e-17	$cmodel
C834	VDD#296	VSS	5.94258e-17	$cmodel
C835	BL<32>#3	VSS	4.79226e-17	$cmodel
C836	BL<31>#3	VSS	8.82729e-17	$cmodel
C837	VDD#286	VSS	2.49053e-17	$cmodel
C838	VDD#287	VSS	2.50001e-17	$cmodel
C839	BLB<31>#3	VSS	1.28016e-16	$cmodel
C840	BLB<30>#2	VSS	7.41074e-17	$cmodel
C841	VDD#277	VSS	5.91314e-17	$cmodel
C842	VDD#278	VSS	5.94258e-17	$cmodel
C843	BL<30>#3	VSS	4.79226e-17	$cmodel
C844	BL<29>#3	VSS	8.82729e-17	$cmodel
C845	VDD#268	VSS	2.49053e-17	$cmodel
C846	VDD#269	VSS	2.50001e-17	$cmodel
C847	BLB<29>#3	VSS	1.28016e-16	$cmodel
C848	BLB<28>#2	VSS	7.41074e-17	$cmodel
C849	VDD#259	VSS	5.91314e-17	$cmodel
C850	VDD#260	VSS	5.94258e-17	$cmodel
C851	BL<28>#3	VSS	4.79226e-17	$cmodel
C852	BL<27>#3	VSS	8.82729e-17	$cmodel
C853	VDD#250	VSS	2.49053e-17	$cmodel
C854	VDD#251	VSS	2.50001e-17	$cmodel
C855	BLB<27>#3	VSS	1.28016e-16	$cmodel
C856	BLB<26>#2	VSS	7.41074e-17	$cmodel
C857	VDD#241	VSS	5.91314e-17	$cmodel
C858	VDD#242	VSS	5.94258e-17	$cmodel
C859	BL<26>#3	VSS	4.79226e-17	$cmodel
C860	BL<25>#3	VSS	8.82729e-17	$cmodel
C861	VDD#232	VSS	2.49053e-17	$cmodel
C862	VDD#233	VSS	2.50001e-17	$cmodel
C863	BLB<25>#3	VSS	1.28016e-16	$cmodel
C864	BLB<24>#2	VSS	7.41074e-17	$cmodel
C865	VDD#223	VSS	5.91314e-17	$cmodel
C866	VDD#224	VSS	5.94258e-17	$cmodel
C867	BL<24>#3	VSS	4.79226e-17	$cmodel
C868	BL<23>#3	VSS	8.82729e-17	$cmodel
C869	VDD#214	VSS	2.49053e-17	$cmodel
C870	VDD#215	VSS	2.50001e-17	$cmodel
C871	BLB<23>#3	VSS	1.28016e-16	$cmodel
C872	BLB<22>#2	VSS	7.41074e-17	$cmodel
C873	VDD#205	VSS	5.91314e-17	$cmodel
C874	VDD#206	VSS	5.94258e-17	$cmodel
C875	BL<22>#3	VSS	4.79226e-17	$cmodel
C876	BL<21>#3	VSS	8.82729e-17	$cmodel
C877	VDD#196	VSS	2.49053e-17	$cmodel
C878	VDD#197	VSS	2.50001e-17	$cmodel
C879	BLB<21>#3	VSS	1.28016e-16	$cmodel
C880	BLB<20>#2	VSS	7.41074e-17	$cmodel
C881	VDD#187	VSS	5.91314e-17	$cmodel
C882	VDD#188	VSS	5.94258e-17	$cmodel
C883	BL<20>#3	VSS	4.79226e-17	$cmodel
C884	BL<19>#3	VSS	8.82729e-17	$cmodel
C885	VDD#178	VSS	2.49053e-17	$cmodel
C886	VDD#179	VSS	2.50001e-17	$cmodel
C887	BLB<19>#3	VSS	1.28016e-16	$cmodel
C888	BLB<18>#2	VSS	7.41074e-17	$cmodel
C889	VDD#169	VSS	5.91314e-17	$cmodel
C890	VDD#170	VSS	5.94258e-17	$cmodel
C891	BL<18>#3	VSS	4.79226e-17	$cmodel
C892	BL<17>#3	VSS	8.82729e-17	$cmodel
C893	VDD#160	VSS	2.49053e-17	$cmodel
C894	VDD#161	VSS	2.50001e-17	$cmodel
C895	BLB<17>#3	VSS	1.28016e-16	$cmodel
C896	BLB<16>#2	VSS	7.41074e-17	$cmodel
C897	VDD#151	VSS	5.91314e-17	$cmodel
C898	VDD#152	VSS	5.94258e-17	$cmodel
C899	BL<16>#3	VSS	4.79226e-17	$cmodel
C900	BL<15>#3	VSS	8.82729e-17	$cmodel
C901	VDD#142	VSS	2.49053e-17	$cmodel
C902	VDD#143	VSS	2.50001e-17	$cmodel
C903	BLB<15>#3	VSS	1.28016e-16	$cmodel
C904	BLB<14>#2	VSS	7.41074e-17	$cmodel
C905	VDD#133	VSS	5.91314e-17	$cmodel
C906	VDD#134	VSS	5.94258e-17	$cmodel
C907	BL<14>#3	VSS	4.79226e-17	$cmodel
C908	BL<13>#3	VSS	8.82729e-17	$cmodel
C909	VDD#124	VSS	2.49053e-17	$cmodel
C910	VDD#125	VSS	2.50001e-17	$cmodel
C911	BLB<13>#3	VSS	1.28016e-16	$cmodel
C912	BLB<12>#2	VSS	7.41074e-17	$cmodel
C913	VDD#115	VSS	5.91314e-17	$cmodel
C914	VDD#116	VSS	5.94258e-17	$cmodel
C915	BL<12>#3	VSS	4.79226e-17	$cmodel
C916	BL<11>#3	VSS	8.82729e-17	$cmodel
C917	VDD#106	VSS	2.49053e-17	$cmodel
C918	VDD#107	VSS	2.50001e-17	$cmodel
C919	BLB<11>#3	VSS	1.28016e-16	$cmodel
C920	BLB<10>#2	VSS	7.41074e-17	$cmodel
C921	VDD#97	VSS	5.91314e-17	$cmodel
C922	VDD#98	VSS	5.94258e-17	$cmodel
C923	BL<10>#3	VSS	4.79226e-17	$cmodel
C924	BL<9>#3	VSS	8.82729e-17	$cmodel
C925	VDD#88	VSS	2.49053e-17	$cmodel
C926	VDD#89	VSS	2.50001e-17	$cmodel
C927	BLB<9>#3	VSS	1.28016e-16	$cmodel
C928	BLB<8>#2	VSS	7.41074e-17	$cmodel
C929	VDD#79	VSS	5.91314e-17	$cmodel
C930	VDD#80	VSS	5.94258e-17	$cmodel
C931	BL<8>#3	VSS	4.79226e-17	$cmodel
C932	BL<7>#3	VSS	8.82729e-17	$cmodel
C933	VDD#70	VSS	2.49053e-17	$cmodel
C934	VDD#71	VSS	2.50001e-17	$cmodel
C935	BLB<7>#3	VSS	1.28016e-16	$cmodel
C936	BLB<6>#2	VSS	7.41074e-17	$cmodel
C937	VDD#61	VSS	5.91314e-17	$cmodel
C938	VDD#62	VSS	5.94258e-17	$cmodel
C939	BL<6>#3	VSS	4.79226e-17	$cmodel
C940	BL<5>#3	VSS	8.82729e-17	$cmodel
C941	VDD#52	VSS	2.49053e-17	$cmodel
C942	VDD#53	VSS	2.50001e-17	$cmodel
C943	BLB<5>#3	VSS	1.28016e-16	$cmodel
C944	BLB<4>#2	VSS	7.41074e-17	$cmodel
C945	VDD#43	VSS	5.91314e-17	$cmodel
C946	VDD#44	VSS	5.94258e-17	$cmodel
C947	BL<4>#3	VSS	4.79226e-17	$cmodel
C948	BL<3>#3	VSS	8.82729e-17	$cmodel
C949	VDD#34	VSS	2.49053e-17	$cmodel
C950	VDD#35	VSS	2.50001e-17	$cmodel
C951	BLB<3>#3	VSS	1.28016e-16	$cmodel
C952	BLB<2>#2	VSS	7.41074e-17	$cmodel
C953	VDD#25	VSS	5.91314e-17	$cmodel
C954	VDD#26	VSS	5.94258e-17	$cmodel
C955	BL<2>#3	VSS	4.79226e-17	$cmodel
C956	BL<1>#3	VSS	8.82729e-17	$cmodel
C957	VDD#16	VSS	2.49053e-17	$cmodel
C958	VDD#17	VSS	2.50001e-17	$cmodel
C959	BLB<1>#3	VSS	1.28016e-16	$cmodel
C960	BLB<0>#2	VSS	7.41074e-17	$cmodel
C961	VDD#7	VSS	5.92366e-17	$cmodel
C962	VDD#8	VSS	5.93512e-17	$cmodel
C963	BL<0>#3	VSS	4.76327e-17	$cmodel
C964	WL#258	VSS	4.29265e-17	$cmodel
C965	BL<63>#2	VSS	4.8068e-17	$cmodel
C966	VDD#562	VSS	6.97496e-17	$cmodel
C967	VDD#567	VSS	6.74715e-17	$cmodel
C968	VDD#564	VSS	3.49717e-16	$cmodel
C969	BLB<63>#2	VSS	4.48303e-17	$cmodel
C970	WL#257	VSS	5.18494e-17	$cmodel
C971	BLB<62>#2	VSS	9.83082e-17	$cmodel
C972	VDD#561	VSS	3.43036e-17	$cmodel
C973	VDD#556	VSS	3.28846e-17	$cmodel
C974	VDD#558	VSS	3.38815e-16	$cmodel
C975	BL<62>#2	VSS	8.83111e-17	$cmodel
C976	WL#256	VSS	4.90214e-17	$cmodel
C977	BL<61>#2	VSS	4.81344e-17	$cmodel
C978	VDD#550	VSS	6.96263e-17	$cmodel
C979	VDD#555	VSS	6.74595e-17	$cmodel
C980	VDD#552	VSS	3.38672e-16	$cmodel
C981	BLB<61>#2	VSS	4.48322e-17	$cmodel
C982	WL#253	VSS	5.16537e-17	$cmodel
C983	BLB<60>#1	VSS	9.83138e-17	$cmodel
C984	VDD#546	VSS	3.43036e-17	$cmodel
C985	VDD#541	VSS	3.28846e-17	$cmodel
C986	VDD#543	VSS	3.38703e-16	$cmodel
C987	BL<60>#2	VSS	8.83111e-17	$cmodel
C988	WL#249	VSS	4.90214e-17	$cmodel
C989	BL<59>#2	VSS	4.81344e-17	$cmodel
C990	VDD#532	VSS	6.96263e-17	$cmodel
C991	VDD#537	VSS	6.74595e-17	$cmodel
C992	VDD#534	VSS	3.38672e-16	$cmodel
C993	BLB<59>#2	VSS	4.48322e-17	$cmodel
C994	WL#245	VSS	5.16537e-17	$cmodel
C995	BLB<58>#1	VSS	9.83138e-17	$cmodel
C996	VDD#528	VSS	3.43036e-17	$cmodel
C997	VDD#523	VSS	3.28846e-17	$cmodel
C998	VDD#525	VSS	3.38703e-16	$cmodel
C999	BL<58>#2	VSS	8.83111e-17	$cmodel
C1000	WL#241	VSS	4.90214e-17	$cmodel
C1001	BL<57>#2	VSS	4.81344e-17	$cmodel
C1002	VDD#514	VSS	6.96263e-17	$cmodel
C1003	VDD#519	VSS	6.74595e-17	$cmodel
C1004	VDD#516	VSS	3.38672e-16	$cmodel
C1005	BLB<57>#2	VSS	4.48322e-17	$cmodel
C1006	WL#237	VSS	5.16537e-17	$cmodel
C1007	BLB<56>#1	VSS	9.83138e-17	$cmodel
C1008	VDD#510	VSS	3.43036e-17	$cmodel
C1009	VDD#505	VSS	3.28846e-17	$cmodel
C1010	VDD#507	VSS	3.38703e-16	$cmodel
C1011	BL<56>#2	VSS	8.83111e-17	$cmodel
C1012	WL#233	VSS	4.90214e-17	$cmodel
C1013	BL<55>#2	VSS	4.81344e-17	$cmodel
C1014	VDD#496	VSS	6.96263e-17	$cmodel
C1015	VDD#501	VSS	6.74595e-17	$cmodel
C1016	VDD#498	VSS	3.38672e-16	$cmodel
C1017	BLB<55>#2	VSS	4.48322e-17	$cmodel
C1018	WL#229	VSS	5.16537e-17	$cmodel
C1019	BLB<54>#1	VSS	9.83138e-17	$cmodel
C1020	VDD#492	VSS	3.43036e-17	$cmodel
C1021	VDD#487	VSS	3.28846e-17	$cmodel
C1022	VDD#489	VSS	3.38703e-16	$cmodel
C1023	BL<54>#2	VSS	8.83111e-17	$cmodel
C1024	WL#225	VSS	4.90214e-17	$cmodel
C1025	BL<53>#2	VSS	4.81344e-17	$cmodel
C1026	VDD#478	VSS	6.96263e-17	$cmodel
C1027	VDD#483	VSS	6.74595e-17	$cmodel
C1028	VDD#480	VSS	3.38672e-16	$cmodel
C1029	BLB<53>#2	VSS	4.48322e-17	$cmodel
C1030	WL#221	VSS	5.16537e-17	$cmodel
C1031	BLB<52>#1	VSS	9.83138e-17	$cmodel
C1032	VDD#474	VSS	3.43036e-17	$cmodel
C1033	VDD#469	VSS	3.28846e-17	$cmodel
C1034	VDD#471	VSS	3.38703e-16	$cmodel
C1035	BL<52>#2	VSS	8.83111e-17	$cmodel
C1036	WL#217	VSS	4.90214e-17	$cmodel
C1037	BL<51>#2	VSS	4.81344e-17	$cmodel
C1038	VDD#460	VSS	6.96263e-17	$cmodel
C1039	VDD#465	VSS	6.74595e-17	$cmodel
C1040	VDD#462	VSS	3.38672e-16	$cmodel
C1041	BLB<51>#2	VSS	4.48322e-17	$cmodel
C1042	WL#213	VSS	5.16537e-17	$cmodel
C1043	BLB<50>#1	VSS	9.83138e-17	$cmodel
C1044	VDD#456	VSS	3.43036e-17	$cmodel
C1045	VDD#451	VSS	3.28846e-17	$cmodel
C1046	VDD#453	VSS	3.38703e-16	$cmodel
C1047	BL<50>#2	VSS	8.83111e-17	$cmodel
C1048	WL#209	VSS	4.90214e-17	$cmodel
C1049	BL<49>#2	VSS	4.81344e-17	$cmodel
C1050	VDD#442	VSS	6.96263e-17	$cmodel
C1051	VDD#447	VSS	6.74595e-17	$cmodel
C1052	VDD#444	VSS	3.38672e-16	$cmodel
C1053	BLB<49>#2	VSS	4.48322e-17	$cmodel
C1054	WL#205	VSS	5.16537e-17	$cmodel
C1055	BLB<48>#1	VSS	9.83138e-17	$cmodel
C1056	VDD#438	VSS	3.43036e-17	$cmodel
C1057	VDD#433	VSS	3.28846e-17	$cmodel
C1058	VDD#435	VSS	3.38703e-16	$cmodel
C1059	BL<48>#2	VSS	8.83111e-17	$cmodel
C1060	WL#201	VSS	4.90214e-17	$cmodel
C1061	BL<47>#2	VSS	4.81344e-17	$cmodel
C1062	VDD#424	VSS	6.96263e-17	$cmodel
C1063	VDD#429	VSS	6.74595e-17	$cmodel
C1064	VDD#426	VSS	3.38672e-16	$cmodel
C1065	BLB<47>#2	VSS	4.48322e-17	$cmodel
C1066	WL#197	VSS	5.16537e-17	$cmodel
C1067	BLB<46>#1	VSS	9.83138e-17	$cmodel
C1068	VDD#420	VSS	3.43036e-17	$cmodel
C1069	VDD#415	VSS	3.28846e-17	$cmodel
C1070	VDD#417	VSS	3.38703e-16	$cmodel
C1071	BL<46>#2	VSS	8.83111e-17	$cmodel
C1072	WL#193	VSS	4.90214e-17	$cmodel
C1073	BL<45>#2	VSS	4.81344e-17	$cmodel
C1074	VDD#406	VSS	6.96263e-17	$cmodel
C1075	VDD#411	VSS	6.74595e-17	$cmodel
C1076	VDD#408	VSS	3.38672e-16	$cmodel
C1077	BLB<45>#2	VSS	4.48322e-17	$cmodel
C1078	WL#189	VSS	5.16537e-17	$cmodel
C1079	BLB<44>#1	VSS	9.83138e-17	$cmodel
C1080	VDD#402	VSS	3.43036e-17	$cmodel
C1081	VDD#397	VSS	3.28846e-17	$cmodel
C1082	VDD#399	VSS	3.38703e-16	$cmodel
C1083	BL<44>#2	VSS	8.83111e-17	$cmodel
C1084	WL#185	VSS	4.90214e-17	$cmodel
C1085	BL<43>#2	VSS	4.81344e-17	$cmodel
C1086	VDD#388	VSS	6.96263e-17	$cmodel
C1087	VDD#393	VSS	6.74595e-17	$cmodel
C1088	VDD#390	VSS	3.38672e-16	$cmodel
C1089	BLB<43>#2	VSS	4.48322e-17	$cmodel
C1090	WL#181	VSS	5.16537e-17	$cmodel
C1091	BLB<42>#1	VSS	9.83138e-17	$cmodel
C1092	VDD#384	VSS	3.43036e-17	$cmodel
C1093	VDD#379	VSS	3.28846e-17	$cmodel
C1094	VDD#381	VSS	3.38703e-16	$cmodel
C1095	BL<42>#2	VSS	8.83111e-17	$cmodel
C1096	WL#177	VSS	4.90214e-17	$cmodel
C1097	BL<41>#2	VSS	4.81344e-17	$cmodel
C1098	VDD#370	VSS	6.96263e-17	$cmodel
C1099	VDD#375	VSS	6.74595e-17	$cmodel
C1100	VDD#372	VSS	3.38672e-16	$cmodel
C1101	BLB<41>#2	VSS	4.48322e-17	$cmodel
C1102	WL#173	VSS	5.16537e-17	$cmodel
C1103	BLB<40>#1	VSS	9.83138e-17	$cmodel
C1104	VDD#366	VSS	3.43036e-17	$cmodel
C1105	VDD#361	VSS	3.28846e-17	$cmodel
C1106	VDD#363	VSS	3.38703e-16	$cmodel
C1107	BL<40>#2	VSS	8.83111e-17	$cmodel
C1108	WL#169	VSS	4.90214e-17	$cmodel
C1109	BL<39>#2	VSS	4.81344e-17	$cmodel
C1110	VDD#352	VSS	6.96263e-17	$cmodel
C1111	VDD#357	VSS	6.74595e-17	$cmodel
C1112	VDD#354	VSS	3.38672e-16	$cmodel
C1113	BLB<39>#2	VSS	4.48322e-17	$cmodel
C1114	WL#165	VSS	5.16537e-17	$cmodel
C1115	BLB<38>#1	VSS	9.83138e-17	$cmodel
C1116	VDD#348	VSS	3.43036e-17	$cmodel
C1117	VDD#343	VSS	3.28846e-17	$cmodel
C1118	VDD#345	VSS	3.38703e-16	$cmodel
C1119	BL<38>#2	VSS	8.83111e-17	$cmodel
C1120	WL#161	VSS	4.90214e-17	$cmodel
C1121	BL<37>#2	VSS	4.81344e-17	$cmodel
C1122	VDD#334	VSS	6.96263e-17	$cmodel
C1123	VDD#339	VSS	6.74595e-17	$cmodel
C1124	VDD#336	VSS	3.38672e-16	$cmodel
C1125	BLB<37>#2	VSS	4.48322e-17	$cmodel
C1126	WL#157	VSS	5.16537e-17	$cmodel
C1127	BLB<36>#1	VSS	9.83138e-17	$cmodel
C1128	VDD#330	VSS	3.43036e-17	$cmodel
C1129	VDD#325	VSS	3.28846e-17	$cmodel
C1130	VDD#327	VSS	3.38703e-16	$cmodel
C1131	BL<36>#2	VSS	8.83111e-17	$cmodel
C1132	WL#153	VSS	4.90214e-17	$cmodel
C1133	BL<35>#2	VSS	4.81344e-17	$cmodel
C1134	VDD#316	VSS	6.96263e-17	$cmodel
C1135	VDD#321	VSS	6.74595e-17	$cmodel
C1136	VDD#318	VSS	3.38672e-16	$cmodel
C1137	BLB<35>#2	VSS	4.48322e-17	$cmodel
C1138	WL#149	VSS	5.16537e-17	$cmodel
C1139	BLB<34>#1	VSS	9.83138e-17	$cmodel
C1140	VDD#312	VSS	3.43036e-17	$cmodel
C1141	VDD#307	VSS	3.28846e-17	$cmodel
C1142	VDD#309	VSS	3.38703e-16	$cmodel
C1143	BL<34>#2	VSS	8.83111e-17	$cmodel
C1144	WL#145	VSS	4.90214e-17	$cmodel
C1145	BL<33>#2	VSS	4.81344e-17	$cmodel
C1146	VDD#298	VSS	6.96263e-17	$cmodel
C1147	VDD#303	VSS	6.74595e-17	$cmodel
C1148	VDD#300	VSS	3.38672e-16	$cmodel
C1149	BLB<33>#2	VSS	4.48322e-17	$cmodel
C1150	WL#141	VSS	5.16537e-17	$cmodel
C1151	BLB<32>#1	VSS	9.83138e-17	$cmodel
C1152	VDD#294	VSS	3.43036e-17	$cmodel
C1153	VDD#289	VSS	3.28846e-17	$cmodel
C1154	VDD#291	VSS	3.38704e-16	$cmodel
C1155	BL<32>#2	VSS	8.83111e-17	$cmodel
C1156	WL#137	VSS	4.90214e-17	$cmodel
C1157	BL<31>#2	VSS	4.81344e-17	$cmodel
C1158	VDD#280	VSS	6.96263e-17	$cmodel
C1159	VDD#285	VSS	6.74595e-17	$cmodel
C1160	VDD#282	VSS	3.38672e-16	$cmodel
C1161	BLB<31>#2	VSS	4.48322e-17	$cmodel
C1162	WL#133	VSS	5.16537e-17	$cmodel
C1163	BLB<30>#1	VSS	9.83138e-17	$cmodel
C1164	VDD#276	VSS	3.43036e-17	$cmodel
C1165	VDD#271	VSS	3.28846e-17	$cmodel
C1166	VDD#273	VSS	3.38703e-16	$cmodel
C1167	BL<30>#2	VSS	8.83111e-17	$cmodel
C1168	WL#129	VSS	4.90214e-17	$cmodel
C1169	BL<29>#2	VSS	4.81344e-17	$cmodel
C1170	VDD#262	VSS	6.96263e-17	$cmodel
C1171	VDD#267	VSS	6.74595e-17	$cmodel
C1172	VDD#264	VSS	3.38672e-16	$cmodel
C1173	BLB<29>#2	VSS	4.48322e-17	$cmodel
C1174	WL#125	VSS	5.16537e-17	$cmodel
C1175	BLB<28>#1	VSS	9.83138e-17	$cmodel
C1176	VDD#258	VSS	3.43036e-17	$cmodel
C1177	VDD#253	VSS	3.28846e-17	$cmodel
C1178	VDD#255	VSS	3.38703e-16	$cmodel
C1179	BL<28>#2	VSS	8.83111e-17	$cmodel
C1180	WL#121	VSS	4.90214e-17	$cmodel
C1181	BL<27>#2	VSS	4.81344e-17	$cmodel
C1182	VDD#244	VSS	6.96263e-17	$cmodel
C1183	VDD#249	VSS	6.74595e-17	$cmodel
C1184	VDD#246	VSS	3.38672e-16	$cmodel
C1185	BLB<27>#2	VSS	4.48322e-17	$cmodel
C1186	WL#117	VSS	5.16537e-17	$cmodel
C1187	BLB<26>#1	VSS	9.83138e-17	$cmodel
C1188	VDD#240	VSS	3.43036e-17	$cmodel
C1189	VDD#235	VSS	3.28846e-17	$cmodel
C1190	VDD#237	VSS	3.38703e-16	$cmodel
C1191	BL<26>#2	VSS	8.83111e-17	$cmodel
C1192	WL#113	VSS	4.90214e-17	$cmodel
C1193	BL<25>#2	VSS	4.81344e-17	$cmodel
C1194	VDD#226	VSS	6.96263e-17	$cmodel
C1195	VDD#231	VSS	6.74595e-17	$cmodel
C1196	VDD#228	VSS	3.38672e-16	$cmodel
C1197	BLB<25>#2	VSS	4.48322e-17	$cmodel
C1198	WL#109	VSS	5.16537e-17	$cmodel
C1199	BLB<24>#1	VSS	9.83138e-17	$cmodel
C1200	VDD#222	VSS	3.43036e-17	$cmodel
C1201	VDD#217	VSS	3.28846e-17	$cmodel
C1202	VDD#219	VSS	3.38703e-16	$cmodel
C1203	BL<24>#2	VSS	8.83111e-17	$cmodel
C1204	WL#105	VSS	4.90214e-17	$cmodel
C1205	BL<23>#2	VSS	4.81344e-17	$cmodel
C1206	VDD#208	VSS	6.96263e-17	$cmodel
C1207	VDD#213	VSS	6.74595e-17	$cmodel
C1208	VDD#210	VSS	3.38672e-16	$cmodel
C1209	BLB<23>#2	VSS	4.48322e-17	$cmodel
C1210	WL#101	VSS	5.16537e-17	$cmodel
C1211	BLB<22>#1	VSS	9.83138e-17	$cmodel
C1212	VDD#204	VSS	3.43036e-17	$cmodel
C1213	VDD#199	VSS	3.28846e-17	$cmodel
C1214	VDD#201	VSS	3.38703e-16	$cmodel
C1215	BL<22>#2	VSS	8.83111e-17	$cmodel
C1216	WL#97	VSS	4.90214e-17	$cmodel
C1217	BL<21>#2	VSS	4.81344e-17	$cmodel
C1218	VDD#190	VSS	6.96263e-17	$cmodel
C1219	VDD#195	VSS	6.74595e-17	$cmodel
C1220	VDD#192	VSS	3.38672e-16	$cmodel
C1221	BLB<21>#2	VSS	4.48322e-17	$cmodel
C1222	WL#93	VSS	5.16537e-17	$cmodel
C1223	BLB<20>#1	VSS	9.83138e-17	$cmodel
C1224	VDD#186	VSS	3.43036e-17	$cmodel
C1225	VDD#181	VSS	3.28846e-17	$cmodel
C1226	VDD#183	VSS	3.38703e-16	$cmodel
C1227	BL<20>#2	VSS	8.83111e-17	$cmodel
C1228	WL#89	VSS	4.90214e-17	$cmodel
C1229	BL<19>#2	VSS	4.81344e-17	$cmodel
C1230	VDD#172	VSS	6.96263e-17	$cmodel
C1231	VDD#177	VSS	6.74595e-17	$cmodel
C1232	VDD#174	VSS	3.38672e-16	$cmodel
C1233	BLB<19>#2	VSS	4.48322e-17	$cmodel
C1234	WL#85	VSS	5.16537e-17	$cmodel
C1235	BLB<18>#1	VSS	9.83138e-17	$cmodel
C1236	VDD#168	VSS	3.43036e-17	$cmodel
C1237	VDD#163	VSS	3.28846e-17	$cmodel
C1238	VDD#165	VSS	3.38703e-16	$cmodel
C1239	BL<18>#2	VSS	8.83111e-17	$cmodel
C1240	WL#81	VSS	4.90214e-17	$cmodel
C1241	BL<17>#2	VSS	4.81344e-17	$cmodel
C1242	VDD#154	VSS	6.96263e-17	$cmodel
C1243	VDD#159	VSS	6.74595e-17	$cmodel
C1244	VDD#156	VSS	3.38672e-16	$cmodel
C1245	BLB<17>#2	VSS	4.48322e-17	$cmodel
C1246	WL#77	VSS	5.16537e-17	$cmodel
C1247	BLB<16>#1	VSS	9.83138e-17	$cmodel
C1248	VDD#150	VSS	3.43036e-17	$cmodel
C1249	VDD#145	VSS	3.28846e-17	$cmodel
C1250	VDD#147	VSS	3.38703e-16	$cmodel
C1251	BL<16>#2	VSS	8.83111e-17	$cmodel
C1252	WL#73	VSS	4.90214e-17	$cmodel
C1253	BL<15>#2	VSS	4.81344e-17	$cmodel
C1254	VDD#136	VSS	6.96263e-17	$cmodel
C1255	VDD#141	VSS	6.74595e-17	$cmodel
C1256	VDD#138	VSS	3.38672e-16	$cmodel
C1257	BLB<15>#2	VSS	4.48322e-17	$cmodel
C1258	WL#69	VSS	5.16537e-17	$cmodel
C1259	BLB<14>#1	VSS	9.83138e-17	$cmodel
C1260	VDD#132	VSS	3.43036e-17	$cmodel
C1261	VDD#127	VSS	3.28846e-17	$cmodel
C1262	VDD#129	VSS	3.38703e-16	$cmodel
C1263	BL<14>#2	VSS	8.83111e-17	$cmodel
C1264	WL#65	VSS	4.90214e-17	$cmodel
C1265	BL<13>#2	VSS	4.81344e-17	$cmodel
C1266	VDD#118	VSS	6.96263e-17	$cmodel
C1267	VDD#123	VSS	6.74595e-17	$cmodel
C1268	VDD#120	VSS	3.38672e-16	$cmodel
C1269	BLB<13>#2	VSS	4.48322e-17	$cmodel
C1270	WL#61	VSS	5.16537e-17	$cmodel
C1271	BLB<12>#1	VSS	9.83138e-17	$cmodel
C1272	VDD#114	VSS	3.43036e-17	$cmodel
C1273	VDD#109	VSS	3.28846e-17	$cmodel
C1274	VDD#111	VSS	3.38703e-16	$cmodel
C1275	BL<12>#2	VSS	8.83111e-17	$cmodel
C1276	WL#57	VSS	4.90214e-17	$cmodel
C1277	BL<11>#2	VSS	4.81344e-17	$cmodel
C1278	VDD#100	VSS	6.96263e-17	$cmodel
C1279	VDD#105	VSS	6.74595e-17	$cmodel
C1280	VDD#102	VSS	3.38672e-16	$cmodel
C1281	BLB<11>#2	VSS	4.48322e-17	$cmodel
C1282	WL#53	VSS	5.16537e-17	$cmodel
C1283	BLB<10>#1	VSS	9.83138e-17	$cmodel
C1284	VDD#96	VSS	3.43036e-17	$cmodel
C1285	VDD#91	VSS	3.28846e-17	$cmodel
C1286	VDD#93	VSS	3.38703e-16	$cmodel
C1287	BL<10>#2	VSS	8.83111e-17	$cmodel
C1288	WL#49	VSS	4.90214e-17	$cmodel
C1289	BL<9>#2	VSS	4.81344e-17	$cmodel
C1290	VDD#82	VSS	6.96263e-17	$cmodel
C1291	VDD#87	VSS	6.74595e-17	$cmodel
C1292	VDD#84	VSS	3.38672e-16	$cmodel
C1293	BLB<9>#2	VSS	4.48322e-17	$cmodel
C1294	WL#45	VSS	5.16537e-17	$cmodel
C1295	BLB<8>#1	VSS	9.83138e-17	$cmodel
C1296	VDD#78	VSS	3.43036e-17	$cmodel
C1297	VDD#73	VSS	3.28846e-17	$cmodel
C1298	VDD#75	VSS	3.38703e-16	$cmodel
C1299	BL<8>#2	VSS	8.83111e-17	$cmodel
C1300	WL#41	VSS	4.90214e-17	$cmodel
C1301	BL<7>#2	VSS	4.81344e-17	$cmodel
C1302	VDD#64	VSS	6.96263e-17	$cmodel
C1303	VDD#69	VSS	6.74595e-17	$cmodel
C1304	VDD#66	VSS	3.38672e-16	$cmodel
C1305	BLB<7>#2	VSS	4.48322e-17	$cmodel
C1306	WL#37	VSS	5.16537e-17	$cmodel
C1307	BLB<6>#1	VSS	9.83138e-17	$cmodel
C1308	VDD#60	VSS	3.43036e-17	$cmodel
C1309	VDD#55	VSS	3.28846e-17	$cmodel
C1310	VDD#57	VSS	3.38703e-16	$cmodel
C1311	BL<6>#2	VSS	8.83111e-17	$cmodel
C1312	WL#33	VSS	4.90214e-17	$cmodel
C1313	BL<5>#2	VSS	4.81344e-17	$cmodel
C1314	VDD#46	VSS	6.96263e-17	$cmodel
C1315	VDD#51	VSS	6.74595e-17	$cmodel
C1316	VDD#48	VSS	3.38672e-16	$cmodel
C1317	BLB<5>#2	VSS	4.48322e-17	$cmodel
C1318	WL#29	VSS	5.16537e-17	$cmodel
C1319	BLB<4>#1	VSS	9.83138e-17	$cmodel
C1320	VDD#42	VSS	3.43036e-17	$cmodel
C1321	VDD#37	VSS	3.28846e-17	$cmodel
C1322	VDD#39	VSS	3.38703e-16	$cmodel
C1323	BL<4>#2	VSS	8.83111e-17	$cmodel
C1324	WL#25	VSS	4.90214e-17	$cmodel
C1325	BL<3>#2	VSS	4.81344e-17	$cmodel
C1326	VDD#28	VSS	6.96263e-17	$cmodel
C1327	VDD#33	VSS	6.74595e-17	$cmodel
C1328	VDD#30	VSS	3.38672e-16	$cmodel
C1329	BLB<3>#2	VSS	4.48322e-17	$cmodel
C1330	WL#21	VSS	5.16537e-17	$cmodel
C1331	BLB<2>#1	VSS	9.83138e-17	$cmodel
C1332	VDD#24	VSS	3.43036e-17	$cmodel
C1333	VDD#19	VSS	3.28846e-17	$cmodel
C1334	VDD#21	VSS	3.38703e-16	$cmodel
C1335	BL<2>#2	VSS	8.83111e-17	$cmodel
C1336	WL#17	VSS	4.90214e-17	$cmodel
C1337	BL<1>#2	VSS	4.81344e-17	$cmodel
C1338	VDD#10	VSS	6.96263e-17	$cmodel
C1339	VDD#15	VSS	6.74595e-17	$cmodel
C1340	VDD#12	VSS	3.38672e-16	$cmodel
C1341	BLB<1>#2	VSS	4.48322e-17	$cmodel
C1342	WL#13	VSS	5.16537e-17	$cmodel
C1343	BLB<0>#1	VSS	9.83138e-17	$cmodel
C1344	VDD#6	VSS	3.43913e-17	$cmodel
C1345	VDD#1	VSS	3.28827e-17	$cmodel
C1346	VDD#3	VSS	3.50866e-16	$cmodel
C1347	BL<0>#2	VSS	8.81323e-17	$cmodel
C1348	WL#9	VSS	1.76204e-16	$cmodel
C1349	VDD#565	VSS	7.19549e-17	$cmodel
C1350	I0<7>/I1<7>/Q#4	VSS	5.63023e-17	$cmodel
C1351	I0<7>/I1<7>/Q#5	VSS	5.15049e-17	$cmodel
C1352	VDD#566	VSS	2.86808e-17	$cmodel
C1353	VDD#563	VSS	2.80432e-17	$cmodel
C1354	I0<7>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1355	I0<7>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1356	I0<7>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1357	VDD#559	VSS	7.04051e-17	$cmodel
C1358	VDD#560	VSS	2.80562e-17	$cmodel
C1359	I0<7>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1360	I0<7>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1361	VDD#557	VSS	2.87131e-17	$cmodel
C1362	I0<7>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1363	I0<7>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1364	VDD#553	VSS	7.18603e-17	$cmodel
C1365	I0<7>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1366	VDD#554	VSS	2.87175e-17	$cmodel
C1367	VDD#551	VSS	2.80432e-17	$cmodel
C1368	I0<7>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1369	I0<7>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1370	I0<7>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1371	VDD#544	VSS	7.02553e-17	$cmodel
C1372	VDD#545	VSS	2.80562e-17	$cmodel
C1373	I0<7>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1374	I0<7>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1375	VDD#542	VSS	2.87131e-17	$cmodel
C1376	I0<7>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1377	I0<7>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1378	VDD#535	VSS	7.18603e-17	$cmodel
C1379	I0<7>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1380	VDD#536	VSS	2.87175e-17	$cmodel
C1381	VDD#533	VSS	2.80432e-17	$cmodel
C1382	I0<7>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1383	I0<7>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1384	I0<7>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1385	VDD#526	VSS	7.02553e-17	$cmodel
C1386	VDD#527	VSS	2.80562e-17	$cmodel
C1387	I0<7>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1388	I0<7>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1389	VDD#524	VSS	2.87131e-17	$cmodel
C1390	I0<7>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1391	I0<7>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1392	VDD#517	VSS	7.18603e-17	$cmodel
C1393	I0<7>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1394	VDD#518	VSS	2.87175e-17	$cmodel
C1395	VDD#515	VSS	2.80432e-17	$cmodel
C1396	I0<7>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1397	I0<7>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1398	I0<7>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1399	VDD#508	VSS	7.02553e-17	$cmodel
C1400	VDD#509	VSS	2.80562e-17	$cmodel
C1401	I0<7>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1402	I0<7>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1403	VDD#506	VSS	2.87131e-17	$cmodel
C1404	I0<7>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1405	I0<6>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1406	VDD#499	VSS	7.18603e-17	$cmodel
C1407	I0<6>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1408	VDD#500	VSS	2.87175e-17	$cmodel
C1409	VDD#497	VSS	2.80432e-17	$cmodel
C1410	I0<6>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1411	I0<6>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1412	I0<6>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1413	VDD#490	VSS	7.02553e-17	$cmodel
C1414	VDD#491	VSS	2.80562e-17	$cmodel
C1415	I0<6>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1416	I0<6>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1417	VDD#488	VSS	2.87131e-17	$cmodel
C1418	I0<6>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1419	I0<6>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1420	VDD#481	VSS	7.18603e-17	$cmodel
C1421	I0<6>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1422	VDD#482	VSS	2.87175e-17	$cmodel
C1423	VDD#479	VSS	2.80432e-17	$cmodel
C1424	I0<6>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1425	I0<6>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1426	I0<6>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1427	VDD#472	VSS	7.02553e-17	$cmodel
C1428	VDD#473	VSS	2.80562e-17	$cmodel
C1429	I0<6>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1430	I0<6>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1431	VDD#470	VSS	2.87131e-17	$cmodel
C1432	I0<6>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1433	I0<6>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1434	VDD#463	VSS	7.18603e-17	$cmodel
C1435	I0<6>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1436	VDD#464	VSS	2.87175e-17	$cmodel
C1437	VDD#461	VSS	2.80432e-17	$cmodel
C1438	I0<6>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1439	I0<6>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1440	I0<6>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1441	VDD#454	VSS	7.02553e-17	$cmodel
C1442	VDD#455	VSS	2.80562e-17	$cmodel
C1443	I0<6>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1444	I0<6>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1445	VDD#452	VSS	2.87131e-17	$cmodel
C1446	I0<6>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1447	I0<6>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1448	VDD#445	VSS	7.18603e-17	$cmodel
C1449	I0<6>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1450	VDD#446	VSS	2.87175e-17	$cmodel
C1451	VDD#443	VSS	2.80432e-17	$cmodel
C1452	I0<6>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1453	I0<6>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1454	I0<6>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1455	VDD#436	VSS	7.02553e-17	$cmodel
C1456	VDD#437	VSS	2.80562e-17	$cmodel
C1457	I0<6>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1458	I0<6>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1459	VDD#434	VSS	2.87131e-17	$cmodel
C1460	I0<6>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1461	I0<5>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1462	VDD#427	VSS	7.18603e-17	$cmodel
C1463	I0<5>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1464	VDD#428	VSS	2.87175e-17	$cmodel
C1465	VDD#425	VSS	2.80432e-17	$cmodel
C1466	I0<5>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1467	I0<5>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1468	I0<5>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1469	VDD#418	VSS	7.02553e-17	$cmodel
C1470	VDD#419	VSS	2.80562e-17	$cmodel
C1471	I0<5>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1472	I0<5>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1473	VDD#416	VSS	2.87131e-17	$cmodel
C1474	I0<5>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1475	I0<5>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1476	VDD#409	VSS	7.18603e-17	$cmodel
C1477	I0<5>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1478	VDD#410	VSS	2.87175e-17	$cmodel
C1479	VDD#407	VSS	2.80432e-17	$cmodel
C1480	I0<5>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1481	I0<5>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1482	I0<5>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1483	VDD#400	VSS	7.02553e-17	$cmodel
C1484	VDD#401	VSS	2.80562e-17	$cmodel
C1485	I0<5>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1486	I0<5>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1487	VDD#398	VSS	2.87131e-17	$cmodel
C1488	I0<5>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1489	I0<5>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1490	VDD#391	VSS	7.18603e-17	$cmodel
C1491	I0<5>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1492	VDD#392	VSS	2.87175e-17	$cmodel
C1493	VDD#389	VSS	2.80432e-17	$cmodel
C1494	I0<5>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1495	I0<5>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1496	I0<5>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1497	VDD#382	VSS	7.02553e-17	$cmodel
C1498	VDD#383	VSS	2.80562e-17	$cmodel
C1499	I0<5>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1500	I0<5>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1501	VDD#380	VSS	2.87131e-17	$cmodel
C1502	I0<5>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1503	I0<5>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1504	VDD#373	VSS	7.18603e-17	$cmodel
C1505	I0<5>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1506	VDD#374	VSS	2.87175e-17	$cmodel
C1507	VDD#371	VSS	2.80432e-17	$cmodel
C1508	I0<5>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1509	I0<5>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1510	I0<5>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1511	VDD#364	VSS	7.02553e-17	$cmodel
C1512	VDD#365	VSS	2.80562e-17	$cmodel
C1513	I0<5>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1514	I0<5>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1515	VDD#362	VSS	2.87131e-17	$cmodel
C1516	I0<5>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1517	I0<4>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1518	VDD#355	VSS	7.18603e-17	$cmodel
C1519	I0<4>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1520	VDD#356	VSS	2.87175e-17	$cmodel
C1521	VDD#353	VSS	2.80432e-17	$cmodel
C1522	I0<4>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1523	I0<4>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1524	I0<4>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1525	VDD#346	VSS	7.02553e-17	$cmodel
C1526	VDD#347	VSS	2.80562e-17	$cmodel
C1527	I0<4>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1528	I0<4>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1529	VDD#344	VSS	2.87131e-17	$cmodel
C1530	I0<4>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1531	I0<4>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1532	VDD#337	VSS	7.18603e-17	$cmodel
C1533	I0<4>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1534	VDD#338	VSS	2.87175e-17	$cmodel
C1535	VDD#335	VSS	2.80432e-17	$cmodel
C1536	I0<4>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1537	I0<4>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1538	I0<4>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1539	VDD#328	VSS	7.02553e-17	$cmodel
C1540	VDD#329	VSS	2.80562e-17	$cmodel
C1541	I0<4>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1542	I0<4>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1543	VDD#326	VSS	2.87131e-17	$cmodel
C1544	I0<4>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1545	I0<4>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1546	VDD#319	VSS	7.18603e-17	$cmodel
C1547	I0<4>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1548	VDD#320	VSS	2.87175e-17	$cmodel
C1549	VDD#317	VSS	2.80432e-17	$cmodel
C1550	I0<4>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1551	I0<4>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1552	I0<4>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1553	VDD#310	VSS	7.02553e-17	$cmodel
C1554	VDD#311	VSS	2.80562e-17	$cmodel
C1555	I0<4>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1556	I0<4>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1557	VDD#308	VSS	2.87131e-17	$cmodel
C1558	I0<4>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1559	I0<4>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1560	VDD#301	VSS	7.18603e-17	$cmodel
C1561	I0<4>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1562	VDD#302	VSS	2.87175e-17	$cmodel
C1563	VDD#299	VSS	2.80432e-17	$cmodel
C1564	I0<4>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1565	I0<4>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1566	I0<4>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1567	VDD#292	VSS	7.02553e-17	$cmodel
C1568	VDD#293	VSS	2.80562e-17	$cmodel
C1569	I0<4>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1570	I0<4>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1571	VDD#290	VSS	2.87131e-17	$cmodel
C1572	I0<4>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1573	I0<3>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1574	VDD#283	VSS	7.18603e-17	$cmodel
C1575	I0<3>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1576	VDD#284	VSS	2.87175e-17	$cmodel
C1577	VDD#281	VSS	2.80432e-17	$cmodel
C1578	I0<3>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1579	I0<3>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1580	I0<3>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1581	VDD#274	VSS	7.02553e-17	$cmodel
C1582	VDD#275	VSS	2.80562e-17	$cmodel
C1583	I0<3>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1584	I0<3>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1585	VDD#272	VSS	2.87131e-17	$cmodel
C1586	I0<3>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1587	I0<3>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1588	VDD#265	VSS	7.18603e-17	$cmodel
C1589	I0<3>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1590	VDD#266	VSS	2.87175e-17	$cmodel
C1591	VDD#263	VSS	2.80432e-17	$cmodel
C1592	I0<3>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1593	I0<3>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1594	I0<3>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1595	VDD#256	VSS	7.02553e-17	$cmodel
C1596	VDD#257	VSS	2.80562e-17	$cmodel
C1597	I0<3>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1598	I0<3>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1599	VDD#254	VSS	2.87131e-17	$cmodel
C1600	I0<3>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1601	I0<3>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1602	VDD#247	VSS	7.18603e-17	$cmodel
C1603	I0<3>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1604	VDD#248	VSS	2.87175e-17	$cmodel
C1605	VDD#245	VSS	2.80432e-17	$cmodel
C1606	I0<3>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1607	I0<3>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1608	I0<3>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1609	VDD#238	VSS	7.02553e-17	$cmodel
C1610	VDD#239	VSS	2.80562e-17	$cmodel
C1611	I0<3>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1612	I0<3>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1613	VDD#236	VSS	2.87131e-17	$cmodel
C1614	I0<3>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1615	I0<3>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1616	VDD#229	VSS	7.18603e-17	$cmodel
C1617	I0<3>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1618	VDD#230	VSS	2.87175e-17	$cmodel
C1619	VDD#227	VSS	2.80432e-17	$cmodel
C1620	I0<3>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1621	I0<3>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1622	I0<3>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1623	VDD#220	VSS	7.02553e-17	$cmodel
C1624	VDD#221	VSS	2.80562e-17	$cmodel
C1625	I0<3>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1626	I0<3>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1627	VDD#218	VSS	2.87131e-17	$cmodel
C1628	I0<3>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1629	I0<2>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1630	VDD#211	VSS	7.18603e-17	$cmodel
C1631	I0<2>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1632	VDD#212	VSS	2.87175e-17	$cmodel
C1633	VDD#209	VSS	2.80432e-17	$cmodel
C1634	I0<2>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1635	I0<2>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1636	I0<2>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1637	VDD#202	VSS	7.02553e-17	$cmodel
C1638	VDD#203	VSS	2.80562e-17	$cmodel
C1639	I0<2>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1640	I0<2>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1641	VDD#200	VSS	2.87131e-17	$cmodel
C1642	I0<2>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1643	I0<2>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1644	VDD#193	VSS	7.18603e-17	$cmodel
C1645	I0<2>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1646	VDD#194	VSS	2.87175e-17	$cmodel
C1647	VDD#191	VSS	2.80432e-17	$cmodel
C1648	I0<2>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1649	I0<2>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1650	I0<2>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1651	VDD#184	VSS	7.02553e-17	$cmodel
C1652	VDD#185	VSS	2.80562e-17	$cmodel
C1653	I0<2>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1654	I0<2>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1655	VDD#182	VSS	2.87131e-17	$cmodel
C1656	I0<2>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1657	I0<2>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1658	VDD#175	VSS	7.18603e-17	$cmodel
C1659	I0<2>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1660	VDD#176	VSS	2.87175e-17	$cmodel
C1661	VDD#173	VSS	2.80432e-17	$cmodel
C1662	I0<2>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1663	I0<2>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1664	I0<2>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1665	VDD#166	VSS	7.02553e-17	$cmodel
C1666	VDD#167	VSS	2.80562e-17	$cmodel
C1667	I0<2>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1668	I0<2>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1669	VDD#164	VSS	2.87131e-17	$cmodel
C1670	I0<2>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1671	I0<2>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1672	VDD#157	VSS	7.18603e-17	$cmodel
C1673	I0<2>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1674	VDD#158	VSS	2.87175e-17	$cmodel
C1675	VDD#155	VSS	2.80432e-17	$cmodel
C1676	I0<2>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1677	I0<2>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1678	I0<2>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1679	VDD#148	VSS	7.02553e-17	$cmodel
C1680	VDD#149	VSS	2.80562e-17	$cmodel
C1681	I0<2>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1682	I0<2>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1683	VDD#146	VSS	2.87131e-17	$cmodel
C1684	I0<2>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1685	I0<1>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1686	VDD#139	VSS	7.18603e-17	$cmodel
C1687	I0<1>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1688	VDD#140	VSS	2.87175e-17	$cmodel
C1689	VDD#137	VSS	2.80432e-17	$cmodel
C1690	I0<1>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1691	I0<1>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1692	I0<1>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1693	VDD#130	VSS	7.02553e-17	$cmodel
C1694	VDD#131	VSS	2.80562e-17	$cmodel
C1695	I0<1>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1696	I0<1>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1697	VDD#128	VSS	2.87131e-17	$cmodel
C1698	I0<1>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1699	I0<1>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1700	VDD#121	VSS	7.18603e-17	$cmodel
C1701	I0<1>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1702	VDD#122	VSS	2.87175e-17	$cmodel
C1703	VDD#119	VSS	2.80432e-17	$cmodel
C1704	I0<1>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1705	I0<1>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1706	I0<1>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1707	VDD#112	VSS	7.02553e-17	$cmodel
C1708	VDD#113	VSS	2.80562e-17	$cmodel
C1709	I0<1>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1710	I0<1>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1711	VDD#110	VSS	2.87131e-17	$cmodel
C1712	I0<1>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1713	I0<1>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1714	VDD#103	VSS	7.18603e-17	$cmodel
C1715	I0<1>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1716	VDD#104	VSS	2.87175e-17	$cmodel
C1717	VDD#101	VSS	2.80432e-17	$cmodel
C1718	I0<1>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1719	I0<1>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1720	I0<1>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1721	VDD#94	VSS	7.02553e-17	$cmodel
C1722	VDD#95	VSS	2.80562e-17	$cmodel
C1723	I0<1>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1724	I0<1>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1725	VDD#92	VSS	2.87131e-17	$cmodel
C1726	I0<1>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1727	I0<1>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1728	VDD#85	VSS	7.18603e-17	$cmodel
C1729	I0<1>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1730	VDD#86	VSS	2.87175e-17	$cmodel
C1731	VDD#83	VSS	2.80432e-17	$cmodel
C1732	I0<1>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1733	I0<1>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1734	I0<1>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1735	VDD#76	VSS	7.02553e-17	$cmodel
C1736	VDD#77	VSS	2.80562e-17	$cmodel
C1737	I0<1>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1738	I0<1>/I1<0>/Q#4	VSS	5.14262e-17	$cmodel
C1739	VDD#74	VSS	2.87131e-17	$cmodel
C1740	I0<1>/I1<0>/Q#6	VSS	5.98945e-17	$cmodel
C1741	I0<0>/I1<7>/Q#4	VSS	5.83319e-17	$cmodel
C1742	VDD#67	VSS	7.18603e-17	$cmodel
C1743	I0<0>/I1<7>/Q#5	VSS	5.14966e-17	$cmodel
C1744	VDD#68	VSS	2.87175e-17	$cmodel
C1745	VDD#65	VSS	2.80432e-17	$cmodel
C1746	I0<0>/I1<7>/QB#4	VSS	5.34662e-17	$cmodel
C1747	I0<0>/I1<7>/QB#6	VSS	6.16901e-17	$cmodel
C1748	I0<0>/I1<5>/QB#4	VSS	6.08254e-17	$cmodel
C1749	VDD#58	VSS	7.02553e-17	$cmodel
C1750	VDD#59	VSS	2.80562e-17	$cmodel
C1751	I0<0>/I1<5>/QB#5	VSS	5.29981e-17	$cmodel
C1752	I0<0>/I1<5>/Q#4	VSS	5.14262e-17	$cmodel
C1753	VDD#56	VSS	2.87131e-17	$cmodel
C1754	I0<0>/I1<5>/Q#6	VSS	5.98945e-17	$cmodel
C1755	I0<0>/I1<6>/Q#4	VSS	5.83319e-17	$cmodel
C1756	VDD#49	VSS	7.18603e-17	$cmodel
C1757	I0<0>/I1<6>/Q#5	VSS	5.14966e-17	$cmodel
C1758	VDD#50	VSS	2.87175e-17	$cmodel
C1759	VDD#47	VSS	2.80432e-17	$cmodel
C1760	I0<0>/I1<6>/QB#4	VSS	5.34662e-17	$cmodel
C1761	I0<0>/I1<6>/QB#6	VSS	6.16901e-17	$cmodel
C1762	I0<0>/I1<3>/QB#4	VSS	6.08254e-17	$cmodel
C1763	VDD#40	VSS	7.02553e-17	$cmodel
C1764	VDD#41	VSS	2.80562e-17	$cmodel
C1765	I0<0>/I1<3>/QB#5	VSS	5.29981e-17	$cmodel
C1766	I0<0>/I1<3>/Q#4	VSS	5.14262e-17	$cmodel
C1767	VDD#38	VSS	2.87131e-17	$cmodel
C1768	I0<0>/I1<3>/Q#6	VSS	5.98945e-17	$cmodel
C1769	I0<0>/I1<4>/Q#4	VSS	5.83319e-17	$cmodel
C1770	VDD#31	VSS	7.18603e-17	$cmodel
C1771	I0<0>/I1<4>/Q#5	VSS	5.14966e-17	$cmodel
C1772	VDD#32	VSS	2.87175e-17	$cmodel
C1773	VDD#29	VSS	2.80432e-17	$cmodel
C1774	I0<0>/I1<4>/QB#4	VSS	5.34662e-17	$cmodel
C1775	I0<0>/I1<4>/QB#6	VSS	6.16901e-17	$cmodel
C1776	I0<0>/I1<1>/QB#4	VSS	6.08254e-17	$cmodel
C1777	VDD#22	VSS	7.02553e-17	$cmodel
C1778	VDD#23	VSS	2.80562e-17	$cmodel
C1779	I0<0>/I1<1>/QB#5	VSS	5.29981e-17	$cmodel
C1780	I0<0>/I1<1>/Q#4	VSS	5.14262e-17	$cmodel
C1781	VDD#20	VSS	2.87131e-17	$cmodel
C1782	I0<0>/I1<1>/Q#6	VSS	5.98945e-17	$cmodel
C1783	I0<0>/I1<2>/Q#4	VSS	5.83319e-17	$cmodel
C1784	VDD#13	VSS	7.18603e-17	$cmodel
C1785	I0<0>/I1<2>/Q#5	VSS	5.14966e-17	$cmodel
C1786	VDD#14	VSS	2.87175e-17	$cmodel
C1787	VDD#11	VSS	2.80432e-17	$cmodel
C1788	I0<0>/I1<2>/QB#4	VSS	5.34662e-17	$cmodel
C1789	I0<0>/I1<2>/QB#6	VSS	6.16901e-17	$cmodel
C1790	I0<0>/I1<0>/QB#4	VSS	6.08254e-17	$cmodel
C1791	VDD#4	VSS	7.02424e-17	$cmodel
C1792	VDD#5	VSS	2.80562e-17	$cmodel
C1793	I0<0>/I1<0>/QB#5	VSS	5.29981e-17	$cmodel
C1794	I0<0>/I1<0>/Q#4	VSS	5.13415e-17	$cmodel
C1795	VDD#2	VSS	2.86766e-17	$cmodel
C1796	I0<0>/I1<0>/Q#6	VSS	5.89683e-17	$cmodel
C1797	WL#259	VSS	2.26072e-16	$cmodel
C1798	WL#260	VSS	2.32109e-16	$cmodel
C1799	WL#261	VSS	2.26072e-16	$cmodel
C1800	WL#262	VSS	2.32109e-16	$cmodel
C1801	WL#263	VSS	2.26072e-16	$cmodel
C1802	WL#264	VSS	2.32109e-16	$cmodel
C1803	WL#265	VSS	2.26072e-16	$cmodel
C1804	WL#266	VSS	2.32109e-16	$cmodel
C1805	WL#267	VSS	2.26072e-16	$cmodel
C1806	WL#268	VSS	2.32109e-16	$cmodel
C1807	WL#269	VSS	2.26072e-16	$cmodel
C1808	WL#270	VSS	2.32109e-16	$cmodel
C1809	WL#271	VSS	2.26072e-16	$cmodel
C1810	WL#272	VSS	2.32109e-16	$cmodel
C1811	WL#273	VSS	2.26072e-16	$cmodel
C1812	WL#274	VSS	2.32109e-16	$cmodel
C1813	WL#275	VSS	2.26072e-16	$cmodel
C1814	WL#276	VSS	2.32109e-16	$cmodel
C1815	WL#277	VSS	2.26072e-16	$cmodel
C1816	WL#278	VSS	2.32109e-16	$cmodel
C1817	WL#279	VSS	2.26072e-16	$cmodel
C1818	WL#280	VSS	2.32109e-16	$cmodel
C1819	WL#281	VSS	2.26072e-16	$cmodel
C1820	WL#282	VSS	2.32109e-16	$cmodel
C1821	WL#283	VSS	2.26072e-16	$cmodel
C1822	WL#284	VSS	2.32109e-16	$cmodel
C1823	WL#285	VSS	2.26072e-16	$cmodel
C1824	WL#286	VSS	2.32109e-16	$cmodel
C1825	WL#287	VSS	2.26072e-16	$cmodel
C1826	WL#288	VSS	2.32109e-16	$cmodel
C1827	WL#289	VSS	2.26072e-16	$cmodel
C1828	WL#290	VSS	2.32109e-16	$cmodel
C1829	WL#291	VSS	2.26072e-16	$cmodel
C1830	WL#292	VSS	2.32109e-16	$cmodel
C1831	WL#293	VSS	2.26072e-16	$cmodel
C1832	WL#294	VSS	2.32109e-16	$cmodel
C1833	WL#295	VSS	2.26072e-16	$cmodel
C1834	WL#296	VSS	2.32109e-16	$cmodel
C1835	WL#297	VSS	2.26072e-16	$cmodel
C1836	WL#298	VSS	2.32109e-16	$cmodel
C1837	WL#299	VSS	2.26072e-16	$cmodel
C1838	WL#300	VSS	2.32109e-16	$cmodel
C1839	WL#301	VSS	2.26072e-16	$cmodel
C1840	WL#302	VSS	2.32109e-16	$cmodel
C1841	WL#303	VSS	2.26072e-16	$cmodel
C1842	WL#304	VSS	2.32109e-16	$cmodel
C1843	WL#305	VSS	2.26072e-16	$cmodel
C1844	WL#306	VSS	2.32109e-16	$cmodel
C1845	WL#307	VSS	2.26072e-16	$cmodel
C1846	WL#308	VSS	2.32109e-16	$cmodel
C1847	WL#309	VSS	2.26072e-16	$cmodel
C1848	WL#310	VSS	2.32109e-16	$cmodel
C1849	WL#311	VSS	2.26072e-16	$cmodel
C1850	WL#312	VSS	2.32109e-16	$cmodel
C1851	WL#313	VSS	2.26072e-16	$cmodel
C1852	WL#314	VSS	2.32109e-16	$cmodel
C1853	WL#315	VSS	2.26072e-16	$cmodel
C1854	WL#316	VSS	2.32109e-16	$cmodel
C1855	WL#317	VSS	2.26072e-16	$cmodel
C1856	WL#318	VSS	2.32109e-16	$cmodel
C1857	WL#319	VSS	2.26072e-16	$cmodel
C1858	WL#320	VSS	2.32109e-16	$cmodel
C1859	WL#321	VSS	2.29037e-16	$cmodel
*
*
.ENDS bit_cell_row_64
*
